# ====================================================================
#
#      hal_sh_sh77x9_se77x9.cdl
#
#      Hitachi SE77X9 board HAL package configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  jskov
# Contributors:
# Date:           2001-05-25
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_SH_SH77X9_SE77X9 {
    display       "Hitachi/SH77X9 SE77X9 board"
    parent        CYGPKG_HAL_SH
    requires      ! CYGHWR_HAL_SH_BIGENDIAN
    requires      CYGHWR_HAL_SH_IRQ_USE_IRQLVL
    define_header hal_sh_sh77x9_se77x9.h
    include_dir   cyg/hal
    description   "
        The SE77X9 HAL package provides the support needed to run
        eCos on a Hitachi/SH SE77X9 board."

    compile       hal_diag.c plf_misc.c ser16c550c.c

    implements    CYGINT_HAL_DEBUG_GDB_STUBS
    implements    CYGINT_HAL_DEBUG_GDB_STUBS_BREAK
    implements    CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT
    implements    CYGINT_HAL_VIRTUAL_VECTOR_COMM_BAUD_SUPPORT

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H   <pkgconf/hal_sh.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_sh_sh77x9_se77x9.h>"

        puts $::cdl_header "#define CYGNUM_HAL_SH_SH3_SCIF_PORTS 1"
        puts $::cdl_header "#define CYGHWR_HAL_VSR_TABLE 0x8c000000"
        puts $::cdl_header "#define CYGHWR_HAL_VECTOR_TABLE 0x8c000100"

        puts $::cdl_header "#define HAL_PLATFORM_BOARD  \"SE77X9\""
        puts $::cdl_header "#define HAL_PLATFORM_EXTRA  \"\""
    }

    cdl_option CYGPRI_HAL_SH_SH77X9_VARIANT {
        display       "Board variant"
        flavor        data
        legal_values  {"SE7709RP01" "SE7709SE01" "SE7729SE01"}
        default_value {"SE7709SE01"}
	no_define
	description   "
	    Select the particular board variant used."
    }

    cdl_option CYGPRI_HAL_SH_SH77X9_SUPERIO {
        display       "Board variant has SuperIO controller"
        default_value 0
        compile       smsc37c93x.c
	description   "
	    Set if the board has a SuperIO controller."
    }


    cdl_option CYGPRI_HAL_SH_SH77X9_VARIANT_7709R {
	display       "SE7709RP01 board"
	active_if     { CYGPRI_HAL_SH_SH77X9_VARIANT == "SE7709RP01" }
	calculated    1

	requires      CYGPKG_HAL_SH_7709R
        requires      !CYGPKG_HAL_SH_7709S
        requires      !CYGPKG_HAL_SH_7729
        requires      !CYGPRI_HAL_SH_SH77X9_SUPERIO
        requires      { CYGNUM_HAL_SH_OOC_XTAL_DEFAULT == 20000000 }
	define_proc {
            puts $::cdl_header "#define HAL_PLATFORM_CPU    \"SH 7709R\""
            puts $::cdl_header "#define CYGNUM_HAL_SH_SE77X9_16550_CLOCK 14745000"
            puts $::cdl_header "#define CYGNUM_HAL_SH_SE77X9_16550_BASE 0xb0800000"
            puts $::cdl_header "#define CYGNUM_HAL_SH_SE77X9_LEDS_BASE 0xb1800000"
        }

        description   "Settings for the 7709R variant of the board."
    }

    cdl_option CYGPRI_HAL_SH_SH77X9_VARIANT_7709S {
	display       "SE7709SE01 board"
	active_if     { CYGPRI_HAL_SH_SH77X9_VARIANT == "SE7709SE01" }
	calculated    1
        requires      CYGPRI_HAL_SH_SH77X9_SUPERIO
        requires      !CYGPKG_HAL_SH_7709R
	requires      CYGPKG_HAL_SH_7709S
        requires      !CYGPKG_HAL_SH_7729
	define_proc {
            puts $::cdl_header "#define HAL_PLATFORM_CPU    \"SH 7709S\""
            puts $::cdl_header "#define CYGNUM_HAL_SH_SE77X9_16550_CLOCK 1846200"
            puts $::cdl_header "#define CYGNUM_HAL_SH_SE77X9_16550_BASE 0xb04007f0"
            puts $::cdl_header "#define CYGNUM_HAL_SH_SE77X9_LEDS_BASE 0xb0c00000"
            puts $::cdl_header "#define CYGNUM_HAL_SH_SE77X9_SDRAM_SETUP"
        }

        description   "Settings for the 7709S variant of the board."
    }
	
    cdl_option CYGPRI_HAL_SH_SH77X9_VARIANT_7729 {
	display       "SE7729SE01 board"
	active_if     { CYGPRI_HAL_SH_SH77X9_VARIANT == "SE7729SE01" }
	calculated    1
        requires      CYGPRI_HAL_SH_SH77X9_SUPERIO
        requires      !CYGPKG_HAL_SH_7709R
        requires      !CYGPKG_HAL_SH_7709S
	requires      CYGPKG_HAL_SH_7729
	define_proc {
            puts $::cdl_header "#define HAL_PLATFORM_CPU    \"SH 7729\""
            puts $::cdl_header "#define CYGNUM_HAL_SH_SE77X9_16550_CLOCK 1846200"
            puts $::cdl_header "#define CYGNUM_HAL_SH_SE77X9_16550_BASE 0xb04007f0"
            puts $::cdl_header "#define CYGNUM_HAL_SH_SE77X9_LEDS_BASE 0xb0c00000"
            puts $::cdl_header "#define CYGNUM_HAL_SH_SE77X9_SDRAM_SETUP"
        }

        description   "Settings for the 7729 variant of the board."
    }
	

    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        legal_values  {"RAM" "ROM" "ROMRAM" }
        default_value {"RAM"}
	no_define
	define -file system.h CYG_HAL_STARTUP
        description   "
           When targetting the SE77X9 board it is possible to build
           the system for either RAM bootstrap or ROM bootstrap.
           RAM bootstrap generally requires that the board
           is equipped with ROMs containing a suitable ROM monitor or
           equivalent software that allows GDB to download the eCos
           application on to the board. The ROM bootstrap typically
           requires that the eCos application be blown into EPROMs or
           equivalent technology. ROMRAM bootstrap is similar to ROM
           bootstrap, but everything is copied to RAM before execution 
           starts thus improving performance, but at the cost of an
           increased RAM footprint."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
        display      "Number of communication channels on the board"
        flavor       data
        calculated   2
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
        display          "Debug serial port"
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
           The SE77X9 board has one serial port. This option
           chooses which port will be used to connect to a host
           running GDB."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_DEFAULT {
        display      "Default console channel."
        flavor       data
        calculated   0
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
        display          "Diagnostic serial port"
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_DEFAULT
        description      "
           The SE77X9 board has two serial ports.  This option
           chooses which port will be used for diagnostic output."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CHANNELS_DEFAULT_BAUD {
        display       "Console/GDB serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 57600 115200
        default_value 38400
        define        CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD
        description   "
            This option controls the default baud rate used for the
            Console/GDB connection."
    }

    cdl_component CYGHWR_HAL_SH_PLF_CLOCK_SETTINGS {
        display          "SH on-chip platform clock controls"
        description      "
            The various clocks used by the system are derived from
            these options."
        flavor        none
        no_define
                     
        cdl_option CYGNUM_HAL_SH_OOC_XTAL_DEFAULT {
            display          "SH clock crystal default value"
            flavor           data
            default_value    33333300
            no_define
        }

        cdl_option CYGHWR_HAL_SH_OOC_XTAL {
            display          "SH clock crystal"
            flavor           data
            legal_values     8000000 to 50000000
            default_value    { CYGNUM_HAL_SH_OOC_XTAL_DEFAULT }
            no_define
            description      "
                This option specifies the frequency of the crystal all
                other clocks are derived from."
        }

        cdl_option CYGHWR_HAL_SH_OOC_PLL_1 {
            display          "SH clock PLL circuit 1"
            flavor           data
            default_value    4
            legal_values     { 0 1 2 3 4 6 8 }
            description      "
                This selects the multiplication factor provided by
                PLL1. If PLL1 is disabled via CAP1, this option should
                be set to zero."
        }

        cdl_option CYGHWR_HAL_SH_OOC_PLL_2 {
            display          "SH clock PLL circuit 2"
            flavor           data
            default_value    1
            legal_values     { 0 1 4 }
            no_define
            description      "
                This selects the multiplication factor provided by
                PLL2. If PLL2 is disabled via CAP2, this option should
                be set to zero."
        }

        cdl_option CYGHWR_HAL_SH_OOC_DIVIDER_1 {
            display          "SH clock divider 1"
            flavor           data
            default_value    1
            legal_values     { 1 2 3 4 6 }
            description      "
                This divider option affects the CPU core clock."
        }

        cdl_option CYGHWR_HAL_SH_OOC_DIVIDER_2 {
            display          "SH clock divider 2"
            flavor           data
            default_value    4
            legal_values     { 1 2 3 4 6 }
            description      "
                This divider option affects the peripheral clock."
        }

        cdl_option CYGHWR_HAL_SH_OOC_CLOCK_MODE {
            display          "SH clock mode"
            flavor           data
            default_value    0
            legal_values     { 0 1 2 3 4 7 }
            description      "
                This option must mirror the clock mode hardwired on
                the MD0-MD2 pins of the CPU in order to correctly
                initialize the FRQCR register."
        }
    }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        parent  CYGPKG_NONE
        no_define
        description   "
	    Global build options including control over
	    compiler flags, linker flags and choice of toolchain."


        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "sh-elf" }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { CYGHWR_HAL_SH_BIGENDIAN ? "-mb -m3 -Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -ggdb -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority" : "-ml -m3 -Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -ggdb -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority" }
            description   "
                This option controls the global compiler flags which
                are used to compile all packages by
                default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { CYGHWR_HAL_SH_BIGENDIAN ? "-mb -m3 -ggdb -nostdlib -Wl,--gc-sections -Wl,-static" : "-ml -m3 -ggdb -nostdlib -Wl,--gc-sections -Wl,-static" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }

        cdl_option CYGBLD_BUILD_GDB_STUBS {
            display "Build GDB stub ROM image"
            default_value 0
            requires { CYG_HAL_STARTUP == "ROM" }
            requires CYGSEM_HAL_ROM_MONITOR
            requires CYGBLD_BUILD_COMMON_GDB_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
            requires ! CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT
            requires ! CYGDBG_HAL_DEBUG_GDB_THREAD_SUPPORT
            requires ! CYGDBG_HAL_COMMON_INTERRUPTS_SAVE_MINIMUM_CONTEXT
            requires ! CYGDBG_HAL_COMMON_CONTEXT_SAVE_MINIMUM
            no_define
            description "
                This option enables the building of the GDB stubs for the
                board. The common HAL controls takes care of most of the
                build process, but the final conversion from ELF image to
                binary data is handled by the platform CDL, allowing
                relocation of the data if necessary."

            make -priority 320 {
                <PREFIX>/bin/gdb_module.bin : <PREFIX>/bin/gdb_module.img
                $(OBJCOPY) -O binary $< $@
            }
        }
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { CYG_HAL_STARTUP == "RAM" ? "sh_sh77x9_se77x9_ram" : \
                     CYG_HAL_STARTUP == "ROM" ? "sh_sh77x9_se77x9_rom" : \
                                                "sh_sh77x9_se77x9_romram" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_sh_sh77x9_se77x9_ram.ldi>" : \
                         CYG_HAL_STARTUP == "ROM" ? "<pkgconf/mlt_sh_sh77x9_se77x9_rom.ldi>" : \
                                                    "<pkgconf/mlt_sh_sh77x9_se77x9_romram.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_sh_sh77x9_se77x9_ram.h>" : \
                         CYG_HAL_STARTUP == "ROM" ? "<pkgconf/mlt_sh_sh77x9_se77x9_rom.h>" : \
                                                    "<pkgconf/mlt_sh_sh77x9_se77x9_romram.h>" }
        }
    }

    cdl_option CYGSEM_HAL_USE_ROM_MONITOR {
        display       "Work with a ROM monitor"
        flavor        booldata
        legal_values  { "GDB_stubs" }
        default_value { CYG_HAL_STARTUP == "RAM" ? "GDB_stubs" : 0 }
        requires      { CYG_HAL_STARTUP == "RAM" }
        parent        CYGPKG_HAL_ROM_MONITOR
        description   "
            Support can be enabled for boot ROMs or ROM monitors which contain
            GDB stubs. This support changes various eCos semantics such as
            the encoding of diagnostic output, and the overriding of hardware
            interrupt vectors."
    }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "ROM" }
        description   "
            Enable this option if this program is to be used as a ROM monitor,
            i.e. applications will be loaded into RAM on the board, and this
            ROM monitor may process exceptions or interrupts generated from the
            application. This enables features such as utilizing a separate
            interrupt stack when exceptions are generated."
    }

    cdl_component CYGPKG_REDBOOT_HAL_OPTIONS {
        display       "Redboot HAL options"
        flavor        none
        no_define
        parent        CYGPKG_REDBOOT
        active_if     CYGPKG_REDBOOT
        description   "
            This option lists the target's requirements for a valid Redboot
            configuration."
    
        cdl_option CYGBLD_BUILD_REDBOOT_BIN {
            display       "Build Redboot ROM binary image"
            active_if     CYGBLD_BUILD_REDBOOT
            default_value 1
            no_define
            description "This option enables the conversion of the Redboot ELF
                         image to a binary image suitable for ROM programming."
    
            make -priority 325 {
                <PREFIX>/bin/redboot.bin : <PREFIX>/bin/redboot.elf
                $(OBJCOPY) --strip-debug $< $(@:.bin=.img) 
                $(OBJCOPY) -O srec $< $(@:.bin=.srec)
                $(OBJCOPY) --change-address 0x21000000 -O srec $< $(@:.bin=.eprom.srec)
                $(OBJCOPY) -O binary $< $@
            }
        }
    }
}
