# ====================================================================
#
#      flash_intel_28fxxx.cdl
#
#      FLASH memory - Hardware support for Intel flash parts
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
## Copyright (C) 2002 Gary Thomas
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Contributors:   jskov, gthomas
# Date:           2001-03-21
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_FLASH_INTEL_28FXXX {
    display       "Intel FlashFile FLASH memory support"
    description   "FLASH memory device support for Intel FlashFile"
    parent        CYGPKG_IO_FLASH
    active_if	  CYGPKG_IO_FLASH

    active_if     CYGINT_DEVS_FLASH_INTEL_28FXXX_REQUIRED

    implements    CYGHWR_IO_FLASH_DEVICE

    include_dir   cyg/io

    requires      { CYGINT_DEVS_FLASH_INTEL_VARIANTS != 0 }

    cdl_interface CYGINT_DEVS_FLASH_INTEL_VARIANTS {
        display   "Number of included variants"
    }

    cdl_interface CYGHWR_DEVS_FLASH_INTEL_BUFFERED_WRITES {
        flavor    booldata
        display   "Must support buffered writes"
    }

    cdl_option CYGHWR_DEVS_FLASH_INTEL_28F160S5 {
        display       "Intel 28F160S5 flash memory support"
        default_value 0
        implements    CYGINT_DEVS_FLASH_INTEL_VARIANTS
        implements    CYGHWR_DEVS_FLASH_INTEL_BUFFERED_WRITES
        description   "
            When this option is enabled, the Intel flash driver will be
            able to recognize and handle the 28F160S5
            part in the family."
    }

    cdl_option CYGHWR_DEVS_FLASH_INTEL_28F320B3 {
        display       "Intel 28F320B3 flash memory support"
        default_value 0
        implements    CYGINT_DEVS_FLASH_INTEL_VARIANTS
        description   "
            When this option is enabled, the Intel flash driver will be
            able to recognize and handle the 28F320B3
            part in the family."
    }


    cdl_option CYGHWR_DEVS_FLASH_INTEL_28F320C3 {
        display       "Intel 28F320C3 flash memory support"
        default_value 0
        implements    CYGHWR_IO_FLASH_BLOCK_LOCKING
        implements    CYGINT_DEVS_FLASH_INTEL_VARIANTS
        description   "
            When this option is enabled, the Intel flash driver will be
            able to recognize and handle the 28F320C3
            part in the family."
    }

    cdl_option CYGHWR_DEVS_FLASH_INTEL_28F320S3 {
        display       "Intel 28F320S3 flash memory support"
        default_value 0
        implements    CYGHWR_IO_FLASH_BLOCK_LOCKING
        implements    CYGINT_DEVS_FLASH_INTEL_VARIANTS
        description   "
            When this option is enabled, the Intel flash driver will be
            able to recognize and handle the 28F320S3
            part in the family."
    }
}
