# ====================================================================
#
#      flash_olpcx2294.cdl
#
#      FLASH memory - Hardware support on Olimex LPC-X2294 boards
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2008 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Sergei Gavrikov
# Contributors:   Sergei Gavrikov
# Date:           2008-08-31
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_FLASH_ARM_OLPCX2294 {
    display       "ARM OLPCE2294, OLPCH2294, OLPCL2294 FLASH memory support"

    parent        CYGPKG_IO_FLASH
    active_if     CYGPKG_IO_FLASH
    requires      (CYGPKG_HAL_ARM_LPC2XXX_OLPCE2294 || \
                   CYGPKG_HAL_ARM_LPC2XXX_OLPCH2294 || \
                   CYGPKG_HAL_ARM_LPC2XXX_OLPCL2294)

    compile       arm_olpcx2294_flash.c

    cdl_interface CYGINT_DEVS_FLASH_INTEL_28FXXX_REQUIRED {
        display   "Generic Intel FlashFile driver required"
    }

    implements    CYGINT_DEVS_FLASH_INTEL_28FXXX_REQUIRED

    cdl_option CYGSEM_DEVS_FLASH_INTEL_28F320C3_PARTS {
        display       "Intel 28F320C3 parts used"
        flavor        bool
	calculated    1
        active_if     (CYGPKG_HAL_ARM_LPC2XXX_OLPCE2294 || \
		       CYGPKG_HAL_ARM_LPC2XXX_OLPCH2294)
        requires      CYGHWR_DEVS_FLASH_INTEL_28F320C3
    }

    cdl_option CYGSEM_DEVS_FLASH_INTEL_28F160C3_PARTS {
        display       "Intel 28F160C3 parts used"
        flavor        bool
	calculated    1
        active_if     CYGPKG_HAL_ARM_LPC2XXX_OLPCL2294
        requires      CYGHWR_DEVS_FLASH_INTEL_28F160C3B
    }
}

