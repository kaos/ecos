# ====================================================================
#
#      wallclock.cdl
#
#      eCos wallclock configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  nickg
# Contributors:
# Date:           1999-07-13
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVICES_WALLCLOCK {
    display       "Wallclock device"
    requires      CYGVAR_KERNEL_COUNTERS_CLOCK
    include_dir   cyg/devs
    define_header wallclock.h
    description   "
        The wallclock device provides real time stamps, as opposed
        to the eCos kernel timers which typically just count the
        number of clock ticks since the hardware was powered up.
        Depending on the target platform this device may involve
        interacting with a suitable clock chip, or it may be
        emulated by using the kernel timers."

    cdl_interface CYGINT_WALLCLOCK_IMPLEMENTATIONS {
        display       "Number of wallclock implementations"
        requires      { CYGINT_WALLCLOCK_IMPLEMENTATIONS == 1 }
    }

    cdl_interface CYGINT_WALLCLOCK_HW_IMPLEMENTATIONS {
        display       "Number of hardware wallclock implementations"
    }

    cdl_option CYGIMP_WALLCLOCK_EMULATE {
        display       "Wallclock emulator"
        default_value { CYGINT_WALLCLOCK_HW_IMPLEMENTATIONS == 0 }
        implements    CYGINT_WALLCLOCK_IMPLEMENTATIONS
        compile       emulate.cxx
        description   "
            When this option is enabled, a wallclock device will be
            emulated using the kernel real-time clock."
    }

    cdl_option CYGIMP_WALLCLOCK_SH3 {
        display       "SH3 Wallclock"
        default_value { CYGPKG_HAL_SH }
        active_if     CYGPKG_HAL_SH
        compile       sh3.cxx
        implements    CYGINT_WALLCLOCK_HW_IMPLEMENTATIONS
        implements    CYGINT_WALLCLOCK_IMPLEMENTATIONS
        description   "
            When this option is enabled, a wallclock driver using the
            SH3's on-core Realtime Clock module will be built."
    }


    cdl_component CYGPKG_DEVICES_WALLCLOCK_OPTIONS {
        display "Wallclock build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_DEVICES_WALLCLOCK_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the wallclock device. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_DEVICES_WALLCLOCK_CFLAGS_REMOVE {
            display "Supressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the wallclock device. These flags are removed from
                the set of global flags if present."
        }

        cdl_option CYGPKG_DEVICES_WALLCLOCK_TESTS {
            display "Wallclock tests"
            flavor  data
            no_define
            calculated { "tests/wallclock" }
            description   "
                This option specifies the set of tests for the wallclock device."
        }
    }
}
