# ====================================================================
#
#      serial_h8300.cdl
#
#      eCos serial H8/300 SCI configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Contributors:
# Date:           1999-07-08
#
#####DESCRIPTIONEND####
#
# ====================================================================


cdl_package CYGPKG_IO_SERIAL_H8300_SCI {
    display       "H8/300 SCI serial device drivers"

    parent        CYGPKG_IO_SERIAL_DEVICES
    active_if     CYGPKG_IO_SERIAL
    active_if     CYGPKG_HAL_H8300

    active_if     CYGINT_IO_SERIAL_H8300_SCI_REQUIRED

    requires      CYGPKG_ERROR
    include_dir   cyg/io
    include_files ; # none _exported_ whatsoever
    description   "
           This option enables the serial device drivers for the
           SCI module in Hitachi H8/300 CPUs."
    doc           redirect/ecos-device-drivers.html

    compile       -library=libextras.a h8300_sci_serial.c

    define_proc {
        puts $::cdl_system_header "/***** serial driver proc output start *****/"
        puts $::cdl_system_header "#ifndef CYGDAT_IO_SERIAL_DEVICE_HEADER"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_DEVICE_HEADER <pkgconf/io_serial_h8300_sci.h>"
        puts $::cdl_system_header "#endif"
        puts $::cdl_system_header "/*****  serial driver proc output end  *****/"

        puts $::cdl_header "#include <pkgconf/system.h>";
        puts $::cdl_header "#include CYGDAT_IO_SERIAL_SH_SCI_CFG";
    }

    cdl_component CYGPKG_IO_SERIAL_SH_SCI_OPTIONS {
        display "SCI serial device driver build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."

        cdl_option CYGPKG_IO_SERIAL_SH_SCI_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are
                used in addition to the set of global flags."
        }

        cdl_option CYGPKG_IO_SERIAL_SH_SCI_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are
                removed from the set of global flags if present."
        }
    }
}

# EOF serial_h8300.cdl
