# ====================================================================
#
#      redboot.cdl
#
#      Redboot package configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000, 2001 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Original data:  gthomas
# Contributors:
# Date:           2000-05-01
#
#####DESCRIPTIONEND####
#
# ====================================================================
cdl_package CYGPKG_REDBOOT {
    display       "Redboot ROM monitor"
    define_header redboot.h
    description   "
           This package supports the Redboot \[stand-alone debug monitor\]
           using eCos as the underlying board support mechanism."

    # Since the CYGDAT_REDBOOT_CONSOLE_DEV setting ends up in the platform
    # HAL header, we need to include that here (via hal.h).
    define_proc {
        puts $::cdl_header "#include <pkgconf/hal.h>"
    }

    cdl_component CYGBLD_BUILD_REDBOOT {
        display "Build Redboot ROM ELF image"
        default_value 0
        requires CYGPKG_INFRA
        requires CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
        requires CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT
        requires ! CYGDBG_HAL_DEBUG_GDB_CTRLC_SUPPORT
        requires ! CYGDBG_HAL_COMMON_INTERRUPTS_SAVE_MINIMUM_CONTEXT
        requires ! CYGDBG_HAL_COMMON_CONTEXT_SAVE_MINIMUM

        cdl_option CYGBLD_BUILD_REDBOOT_WITH_THREADS {
            no_define
            active_if { CYG_HAL_STARTUP != "RAM" }
            requires  CYGDBG_HAL_DEBUG_GDB_THREAD_SUPPORT
        }

        no_define
        description "This option enables the building of the Redboot ELF image.
                     The image may require further relocation or symbol
                     stripping before being converted to a binary image.
                     This is handled by a rule in the target CDL."

        compile main.c crc.c
        compile printf.c misc_funs.c io.c parse.c ticks.c xyzModem.c syscall.c
        compile decompress.c
        compile -library=libextras.a load.c 

        make -priority 320 {
            <PREFIX>/bin/redboot.elf : $(PREFIX)/lib/target.ld $(PREFIX)/lib/vectors.o $(PREFIX)/lib/libtarget.a $(PREFIX)/lib/libextras.a
                    @sh -c "mkdir -p $(dir $@)"
                    $(CC) -c $(INCLUDE_PATH) $(CFLAGS) -o $(PREFIX)/lib/version.o $(REPOSITORY)/$(PACKAGE)/src/version.c
	            $(CC) $(LDFLAGS) -L$(PREFIX)/lib -Ttarget.ld -o $@ $(PREFIX)/lib/version.o
        }
    }

    cdl_component CYGPKG_REDBOOT_NETWORKING {
        display       "Build Redboot ROM binary image"
        flavor        bool
        active_if     CYGPKG_IO_ETH_DRIVERS
        default_value 1
	compile net/bootp.c net/udp.c net/ip.c net/pktbuf.c net/cksum.c
	compile net/enet.c net/icmp.c net/tcp.c net/timers.c net/arp.c
	compile net/tftp_client.c net/net_io.c net/inet_addr.c
	compile -library=libextras.a net/ping.c
        description "This option includes networking support in RedBoot."
        define_proc {
            puts $::cdl_system_header "#define CYGNUM_HAL_VIRTUAL_VECTOR_AUX_CHANNELS 1"
        }

        cdl_option CYGNUM_REDBOOT_NETWORKING_TCP_PORT {
            display          "TCP port to listen for incoming connections"
            flavor           data
            default_value    9000
            description      "
               RedBoot will 'listen' on this port for incoming TCP connections.
               This allows outside connections to be made to the platform, either
               for GDB or RedBoot commands."
        }

        cdl_option CYGNUM_REDBOOT_NETWORKING_MAX_PKTBUF {
            display          "Number of \[network\] packet buffers"
            flavor           data
            default_value    4
            legal_values     3 to 8
            description      "
               RedBoot may need to buffer network data to support various connections.
               This option allows control over the number of such buffered packets,
               and in turn, controls the amount of memory used by RedBoot (which
               is not available to user applications).  Each packet buffer takes up
               about 1514 bytes.  Note: there is little need to make this larger
               than the default."
        }
    }

    cdl_option CYGPKG_REDBOOT_ANY_CONSOLE {
        display       "Allow RedBoot to use any I/O channel for it's console."
        flavor        bool
        default_value 1
        description   "
          If this option is enabled then RedBoot will attempt to use all
          defined serial I/O channels for it's console device.  Once input
          arrives at one of these channels then the console will use only
          that port."
    }

    cdl_option CYGPKG_REDBOOT_MAX_CMD_LINE {
        display       "Maximum command line length"
        flavor        data
        default_value 256
        description   "
          This option allows control over how long the CLI command line
          should be.  This space will be allocated statically
          rather than from RedBoot's stack."
    }

    cdl_option CYGNUM_REDBOOT_CLI_IDLE_TIMEOUT {
        display       "Command processing idle timeout (ms)"
        flavor        data
        default_value 10
        description   "
          This option controls the timeout period before the
          command processing is considered 'idle'.  Making this
          number smaller will cause idle processing to take place
          more often, etc.  The default value of 10ms is a reasonable
          tradeoff between responsiveness and overhead."
    }

    cdl_option CYGNUM_REDBOOT_LOAD_ZLIB_BUFFER {
        display       "Size of zlib decompression buffer"
        active_if     CYGPKG_COMPRESS_ZLIB
        flavor        data
        default_value 64
        legal_values  5 to 256
        description   "
            This is the size of the buffer filled with incoming data
            during load before calls are made to the decompressor
            function. For ethernet downloads this can be made bigger
            (at the cost of memory), but for serial downloads on slow
            processors it may be necessary to reduce the size to
            avoid serial overruns. zlib appears to bail out if less than
            five bytes are available initially so this is the minimum."
    }

    cdl_component CYGPKG_REDBOOT_FLASH {
        display       "Allow RedBoot to support FLASH programming"
        flavor        bool
        default_value 1
        active_if     CYGPKG_IO_FLASH
        description   "
          If this option is enabled then RedBoot will provide commands
          to manage images in FLASH memory.  These images can be loaded
          into memory for execution or executed in place."
        compile -library=libextras.a flash.c

        cdl_option CYGBLD_REDBOOT_MIN_IMAGE_SIZE {
            display       "Minimum image size"
            flavor        data
            default_value 0x20000
            description "
              This option controls the minimum length of images kept by
              the FIS.  In particular, it should be large enough to hold
              the RedBoot primary image itself, as well as be a natural
              multiple of the FLASH erase block size."
        }

        cdl_option CYGBLD_REDBOOT_FLASH_BOOT_OFFSET {
            display       "Offset from start of FLASH to RedBoot boot image"
            flavor        data
            default_value CYGNUM_REDBOOT_FLASH_RESERVED_BASE
	    requires      { CYGNUM_REDBOOT_FLASH_RESERVED_BASE <= \
		            CYGBLD_REDBOOT_FLASH_BOOT_OFFSET }
            description "
              This option controls where the RedBoot boot image is located
              relative to the start of FLASH."
        }

        cdl_option CYGNUM_REDBOOT_FLASH_RESERVED_BASE {
            display       "Size of reserved area at start of FLASH"
            flavor        data
            default_value 0
            description "
              This option reserves an area at the start of FLASH where RedBoot
	      will never interfere; it is expected that this area contains
              (non-RedBoot-based) POST code or some other boot monitor that
              executes before RedBoot."
        }

	cdl_component CYGPKG_REDBOOT_FIS_CONTENTS {
	    display       "Flash Image System default directory contents"
	    calculated 1

	    cdl_option CYGOPT_REDBOOT_FIS_RESERVED_BASE {
		display		"Pseudo-file to describe reserved area"
		active_if	{ 0 != CYGNUM_REDBOOT_FLASH_RESERVED_BASE }
		default_value	1
		description "
		    If an area of FLASH is reserved, it is informative to
		    have a fis entry describing it.  This option controls
		    creation of such an entry by default in the fis init
		    command."
	    }

	    cdl_option CYGOPT_REDBOOT_FIS_REDBOOT {
		display		"File to describe RedBoot boot image"
		default_value	1
		description "
		    Normally a ROM-startup RedBoot image is first in the
		    FLASH, and the system boots using that image.  This
		    option controls creation of an entry describing it in
		    the fis init command.  It might be disabled if a
		    platform has an immutable boot image of its own, where
		    we use a POST-startup RedBoot instead, which performs
		    less board initialization."
	    }

	    cdl_component CYGOPT_REDBOOT_FIS_REDBOOT_POST {
		display		"File to describe RedBoot POST-compatible image"
		default_value	!CYGOPT_REDBOOT_FIS_REDBOOT
		description "
		    This option controls creation of an entry describing a
		    POST-startup RedBoot image in the fis init command.
		    Not all platforms support POST-startup.  A platform
		    might have both for testing purposes, where the
		    eventual user would substitute their own POST code for
		    the initial ROM-startup RedBoot, and then jump to the
		    POST-compatible RedBoot immediately following."
		cdl_option CYGNUM_REDBOOT_FIS_REDBOOT_POST_OFFSET {
		    display    "Offset of POST image from FLASH start"
		    flavor     booldata
		    default_value 0
		    requires   { CYGNUM_REDBOOT_FIS_REDBOOT_POST_OFFSET >= \
			         CYGBLD_REDBOOT_FLASH_BOOT_OFFSET }
		    description "
	            This option specifies the offset for a POST image from
		    the start of FLASH.  If unset, then the fis entry
		    describing the POST image will be placed where
		    convenient."
		}
	    }   

	    cdl_option CYGOPT_REDBOOT_FIS_REDBOOT_BACKUP {
		display		"File to describe RedBoot backup image"
		default_value	1
		description "
		    This option controls creation of an entry describing a
		    backup RedBoot image in the fis init command.
		    Conventionally a RAM-startup RedBoot image is kept
		    under this name for use in updating the ROM-based
		    RedBoot that boots the board."
	    }
	}

        cdl_component CYGSEM_REDBOOT_FLASH_CONFIG {
            display       "Keep RedBoot configuration data in FLASH"
            flavor        bool
            default_value 1
            description "
              When this option is enabled, RedBoot will keep configuration
              data in a separate block of FLASH memory.  This data will
              include such items as the node IP address or startup scripts."

            cdl_option CYGNUM_REDBOOT_FLASH_CONFIG_SIZE {
                display       "Length of configuration data in FLASH"
                flavor        data
                default_value 1024
                description "
                  This option is used to control the amount of memory and FLASH
                  to be used for configuration options (persistent storage)."
            }

            cdl_option CYGNUM_REDBOOT_FLASH_SCRIPT_SIZE {
                display       "Length of configuration script(s) in FLASH"
                flavor        data
                default_value 512
                description "
                  This option is used to control the amount of memory and FLASH
                  to be used for configuration options (persistent storage)."
            }
        }

        cdl_option CYGSEM_REDBOOT_FLASH_LOCK_SPECIAL {
            display       "Keep all RedBoot FLASH data blocks locked."
            flavor        bool
            default_value 1
            active_if     { CYGHWR_IO_FLASH_BLOCK_LOCKING != 0 }
            description "
              When this option is enabled, RedBoot will keep configuration
              data and the FIS directory blocks implicitly locked.  While
              this is somewhat safer, it does add overhead during updates."
        }

        cdl_option CYGNUM_REDBOOT_FLASH_SCRIPT_TIMEOUT_RESOLUTION {
            display       "Resolution (in ms) for script timeout value."
            flavor        data
            default_value 1000
            active_if     CYGSEM_REDBOOT_FLASH_CONFIG
            description "
              This option controls the resolution of the script timeout.
              The value is specified in milliseconds (ms), thus to have the
              script timeout be defined in terms of tenths of seconds, use 100."
        }

        cdl_option CYGNUM_REDBOOT_FLASH_SCRIPT_DEFAULT_TIMEOUT {
            display       "Default script timeout value"
            flavor        data
            default_value 10
            active_if     CYGSEM_REDBOOT_FLASH_CONFIG
            description "
              This option is used to set the default timeout for startup
              scripts, when they are enabled."
        }
    }

    cdl_option CYGPRI_REDBOOT_ROM_MONITOR {
        active_if    { CYG_HAL_STARTUP == "ROM" }
        requires     CYGSEM_HAL_ROM_MONITOR
        calculated   1
        no_define
    }

    cdl_option CYGSEM_REDBOOT_BSP_SYSCALLS {
        display       "Allow RedBoot to handle GNUPro application 'syscalls'."
        flavor        bool
        default_value 0
        description   "
          If this option is enabled then RedBoot will install a syscall handler
          to support debugging of applications based on GNUPro newlib/bsp."
    }
}

