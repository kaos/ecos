# ====================================================================
#
#      ser_v85x_v850.cdl
#
#      eCos serial NEC/V850 configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Original data:  gthomas
# Contributors:
# Date:           2000-05-26
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_IO_SERIAL_V85X_V850 {
    display       "NEC V850 serial device drivers"

    parent        CYGPKG_IO_SERIAL_DEVICES
    active_if     CYGPKG_IO_SERIAL
    active_if     CYGPKG_HAL_V85X_V850

    requires      CYGPKG_ERROR
    include_dir   cyg/io
    include_files ; # none _exported_ whatsoever
    description   "
           This option enables the serial device drivers for the
           NEC CEB/V850SA1."
    doc           redirect/ecos-device-drivers.html

    compile       -library=libextras.a   v85x_v850_serial.c

    define_proc {
        puts $::cdl_system_header "/***** serial driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_DEVICE_HEADER <pkgconf/io_serial_v85x_v850.h>"
        puts $::cdl_system_header "/*****  serial driver proc output end  *****/"
    }

    cdl_component CYGPKG_IO_SERIAL_V85X_V850_SERIAL0 {
        display       "NEC V850 serial port 0 driver"
        flavor        bool
        default_value 0
        description   "
            This option includes the serial device driver for the NEC V850
            SA1 (70F3017) and SB1 (70F3033) devices, port 0."
    
        cdl_option CYGDAT_IO_SERIAL_V85X_V850_SERIAL0_NAME {
            display       "Device name for NEC V850 serial port 0 driver"
            flavor        data
            default_value {"\"/dev/ser0\""}
            description   "
                This option specifies the name of the serial device for the 
                NEC V850, port 0."
        }
    
        cdl_option CYGNUM_IO_SERIAL_V85X_V850_SERIAL0_BAUD {
            display       "Baud rate for the NEC V850 serial port 0 driver"
            flavor        data
            legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                          4800 7200 9600 14400 19200 38400 57600 115200
            }
            default_value 38400
            description   "
                This option specifies the default baud rate (speed) for the 
                NEC V850, port 0."
        }
    
        cdl_option CYGNUM_IO_SERIAL_V85X_V850_SERIAL0_BUFSIZE {
            display       "Buffer size for the NEC V850 serial port 0 driver"
            flavor        data
            legal_values  0 to 8192
            default_value 128
            description   "
                This option specifies the size of the internal buffers used 
                for the NEC V850, port 0."
        }
    }

    cdl_component CYGPKG_IO_SERIAL_V85X_V850_TESTING {
        display    "Testing parameters"
        flavor     bool
        calculated 1
        active_if  CYGPKG_IO_SERIAL_V85X_V850_SERIAL0

        cdl_option CYGPRI_SER_TEST_SER_DEV {
            display       "Serial device used for testing"
            flavor        data
            default_value { CYGDAT_IO_SERIAL_V85X_V850_SERIAL0_NAME }
        }

        define_proc {
            puts $::cdl_header "#define CYGPRI_SER_TEST_CRASH_ID \"v85x/v850\""
            puts $::cdl_header "#define CYGPRI_SER_TEST_TTY_DEV  \"/dev/tty0\""
        }
    }

}
