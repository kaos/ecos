# ====================================================================
#
#      i2c.cdl
#
#      Generic I2C package configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 2004 eCosCentric Limited
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):     bartv
# Date:          2004-10-05
#
#####DESCRIPTIONEND####
#========================================================================

cdl_package CYGPKG_IO_I2C {
    display		"I2C support"
    doc			ref/io-i2c.html
    requires		CYGPKG_INFRA CYGPKG_HAL
    hardware
    include_dir		cyg/io
    compile		i2c.cxx
    
    description "
        The generic I2C package provides an API for accessing devices
        attached to an I2C bus. It specifies how I2C bus drivers should
        be written and how I2C devices should be defined. There is also
        support for bit-banged I2C buses."

    cdl_option CYGNUM_I2C_INIT_PRIORITY {
	display		"I2C initialization priority"
	flavor		data
	default_value	{ "CYG_INIT_DRIVERS" }

	description "
            The generic I2C package will initialize each I2C bus during
            system startup, using a prioritized static constructor. This
            option controls the priority that is used. The default value,
            CYG_INIT_DRIVERS, means that I2C buses get initialized early
            on."
    }

    cdl_component CYGPKG_IO_I2C_OPTIONS {
        display "I2C build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building the generic I2C
            package, and details of which tests are built."

        cdl_option CYGPKG_IO_I2C_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the generic I2C package. These flags are
                used in addition to the set of global flags."
        }

        cdl_option CYGPKG_IO_I2C_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the generic I2C package. These flags are
                removed from the set of global flags if present."
        }
    }
}
