# ====================================================================
#
#      ser_arm_integrator.cdl
#
#      eCos serial ARM/INTEGRATOR configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      David A Rusling
# Original data:  David A Rusling
# Contributors:	  Philippe Robin
# Date:           November 7, 2000
#
#####DESCRIPTIONEND####
#
# ====================================================================


cdl_package CYGPKG_IO_SERIAL_ARM_INTEGRATOR {
    display       "ARM INTEGRATOR serial device drivers"

    parent        CYGPKG_IO_SERIAL_DEVICES
    active_if     CYGPKG_IO_SERIAL
    active_if     CYGPKG_HAL_ARM_INTEGRATOR

    requires      CYGPKG_ERROR
    include_dir   cyg/io
    description   "
           This option enables the serial device drivers for the
           ARM INTEGRATOR."
    doc           redirect/ecos-device-drivers.html

    compile       -library=libextras.a   integrator_serial_with_ints.c

    define_proc {
        puts $::cdl_system_header "/***** serial driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_DEVICE_HEADER <pkgconf/io_serial_arm_integrator.h>"
        puts $::cdl_system_header "/*****  serial driver proc output end  *****/"
    }

    cdl_component CYGPKG_IO_SERIAL_ARM_INTEGRATOR_SERIAL0 {
	display       "ARM INTEGRATOR serial port 0 driver"
	flavor        bool
	default_value 1
	description   "
        This option includes the serial device driver for the ARM INTEGRATOR 
        port 0."

	cdl_option CYGDAT_IO_SERIAL_ARM_INTEGRATOR_SERIAL0_NAME {
	    display       "Device name for ARM INTEGRATOR serial port 0 driver"
	    flavor        data
	    default_value {"\"/dev/ser0\""}
	    description   "
            This option specifies the name of the serial device for the 
            ARM INTEGRATOR port 0."
	}

	cdl_option CYGNUM_IO_SERIAL_ARM_INTEGRATOR_SERIAL0_BAUD {
	    display       "Baud rate for the ARM INTEGRATOR serial port 0 driver"
	    flavor        data
	    legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
	    		    4800 7200 9600 14400 19200 38400 57600 115200 234000
			   }
	    default_value 38400
	    description   "
            This option specifies the default baud rate (speed) for the 
            ARM INTEGRATOR port 0."
	}

	cdl_option CYGNUM_IO_SERIAL_ARM_INTEGRATOR_SERIAL0_BUFSIZE {
	    display       "Buffer size for the ARM INTEGRATOR serial port 0 driver"
	    flavor        data
	    legal_values  0 to 8192
	    default_value 128
	    description   "
            This option specifies the size of the internal buffers used 
            for the ARM INTEGRATOR port 0."
	}
    }

    cdl_component CYGPKG_IO_SERIAL_ARM_INTEGRATOR_SERIAL1 {
	display       "ARM INTEGRATOR serial port 1 driver"
	flavor        bool
	default_value 1
	description   "
        This option includes the serial device driver for the ARM INTEGRATOR 
        port 1."

	cdl_option CYGDAT_IO_SERIAL_ARM_INTEGRATOR_SERIAL1_NAME {
	    display       "Device name for ARM INTEGRATOR serial port 1 driver"
	    flavor        data
	    default_value {"\"/dev/ser1\""}
	    description   "
            This option specifies the name of the serial device for the 
            ARM INTEGRATOR port 1."
	}

	cdl_option CYGNUM_IO_SERIAL_ARM_INTEGRATOR_SERIAL1_BAUD {
	    display       "Baud rate for the ARM INTEGRATOR serial port 1 driver"
	    flavor        data
	    legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 234000
            }
	    default_value 38400
	    description   "
            This option specifies the default baud rate (speed) for the
            ARM INTEGRATOR port 1."
	}
    }

    cdl_option CYGNUM_IO_SERIAL_ARM_INTEGRATOR_SERIAL1_BUFSIZE {
        display       "Buffer size for the ARM INTEGRATOR serial port 1 driver"
        flavor        data
        legal_values  0 to 8192
        default_value 128
        description   "
            This option specifies the size of the internal buffers used 
            for the ARM INTEGRATOR port 1."
    }

    cdl_component CYGPKG_IO_SERIAL_ARM_INTEGRATOR_TESTING {
        display    "Testing parameters"
        flavor     bool
        calculated 1
        active_if  CYGPKG_IO_SERIAL_ARM_INTEGRATOR_SERIAL0

# FIXME: I have no idea what the integrator hardware doesn't support -Jifl
#        implements CYGINT_IO_SERIAL_TEST_SKIP_9600
#        implements CYGINT_IO_SERIAL_TEST_SKIP_115200
#        implements CYGINT_IO_SERIAL_TEST_SKIP_PARITY_EVEN
        
        cdl_option CYGPRI_SER_TEST_SER_DEV {
            display       "Serial device used for testing"
            flavor        data
            default_value { CYGDAT_IO_SERIAL_ARM_INTEGRATOR_SERIAL0_NAME }
        }

        define_proc {
            puts $::cdl_header "#define CYGPRI_SER_TEST_CRASH_ID \"arminteg\""
            puts $::cdl_header "#define CYGPRI_SER_TEST_TTY_DEV  \"/dev/tty0\""
        }
    }
}

# EOF ser_arm_integrator.cdl
