# ====================================================================
#
#      hal_mips_tx49.cdl
#
#      MIPS/TX49 variant architectural HAL package configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  bartv, nickg
# Contributors:
# Date:           2000-05-15
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_MIPS_TX49 {
    display       "TX49 variant"
    parent        CYGPKG_HAL_MIPS
    hardware
    include_dir   cyg/hal
    define_header hal_mips_tx49.h
    description   "
           The TX49 architecture HAL package provides generic support
           for this processor architecture. It is also necessary to
           select a specific target platform HAL package."

    cdl_component CYGPKG_HAL_MIPS_TX4955 {
        display       "TX4955 microprocessor"
        default_value 1
        implements    CYGINT_HAL_MIPS_VARIANT
        description "
            The TMPR4955F microprocessor. This is an embedded part that in
            addition to the TX49 processor core has built in peripherals
            such as memory controllers, DMA controllers, serial ports and
            timers/counters."               

        define_proc {
            # Sizes are configurable (on the core). Should be configurable.
            puts $::cdl_header "#define CYGHWR_HAL_DCACHE_SIZE 32768"
            puts $::cdl_header "#define CYGHWR_HAL_ICACHE_SIZE 32768"
        }

        cdl_option CYGHWR_HAL_MIPS_64BIT {
            display    "Variant 64 bit architecture support"
            description "
                While the TX49 is a 64bit CPU, only its 32bit mode is
                currently supported in eCos."
            calculated 0
        }

        # This is optional (on the core). Should be configurable.
        cdl_option CYGHWR_HAL_MIPS_FPU {
            display    "Variant FPU support"
            calculated 1
        }

        cdl_interface CYGINT_HAL_MIPS_FPU_64BIT {
            display "Variant 64 bit FPU support interface"
        }

        cdl_option CYGHWR_HAL_MIPS_FPU_64BIT {
            display    "Variant 64 bit FPU support"
            calculated { CYGINT_HAL_MIPS_FPU_64BIT == 1 ? 1 : 0 }
        }

        cdl_option CYGHWR_HAL_MIPS_FPU_32BIT {
            display    "Variant 32 bit FPU support"
            calculated { CYGINT_HAL_MIPS_FPU_64BIT == 0 ? 1 : 0 }
        }

        # FGRn+1 is most significant part of the FGRn&FGRn+1 pair of FPRn/2
        # This is true for BE mips2 mode at least. Not sure about fp64 mode
        cdl_option CYGPKG_HAL_MIPS_DOUBLE_LSBFIRST {
            active_if CYGHWR_HAL_MIPS_FPU_32BIT
            calculated 1
        }

        cdl_interface CYGINT_HAL_MIPS_MSBFIRST {
            no_define
            display    "CPU Variant big-endian interface"
        }

        cdl_option CYGPKG_HAL_MIPS_MSBFIRST {
            display    "CPU Variant big-endian"
            calculated { CYGINT_HAL_MIPS_MSBFIRST == 0 ? 0 : 1 }
        }

        cdl_option CYGPKG_HAL_MIPS_LSBFIRST {
            display    "CPU Variant little-endian"
            calculated { CYGINT_HAL_MIPS_MSBFIRST != 0 ? 0 : 1 }
        }
    }

    define_proc {
        puts $::cdl_header "#include <pkgconf/hal_mips.h>"
    }

    compile       var_misc.c variant.S

    make {
        <PREFIX>/lib/target.ld: <PACKAGE>/src/mips_tx49.ld
        $(CC) -E -P -Wp,-MD,target.tmp -DEXTRAS=1 -xc $(INCLUDE_PATH) $(CFLAGS) -o $@ $<
        @echo $@ ": \\" > $(notdir $@).deps
        @tail +2 target.tmp >> $(notdir $@).deps
        @echo >> $(notdir $@).deps
        @rm target.tmp
    }

    cdl_option CYGBLD_LINKER_SCRIPT {
        display "Linker script"
        flavor data
	no_define
        calculated  { "src/mips_tx49.ld" }
    }
}
