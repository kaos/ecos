# ====================================================================
#
#      flash_olpcx2294.cdl
#
#      FLASH memory - Hardware support on Olimex LPC-X2294 boards
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
## Copyright (C) 2008 eCosCentric Limited
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Sergei Gavrikov
# Contributors:   Sergei Gavrikov
# Date:           2008-11-28
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_FLASH_ARM_OLPCX2294_V2 {
    display       "Support for FLASH memory parts on OLPC-X2294 boards."

    compile       -library=libextras.a arm_olpcx2294_flash.c

    parent        CYGPKG_IO_FLASH
    active_if     CYGPKG_IO_FLASH

    requires      (CYGPKG_HAL_ARM_LPC2XXX_OLPCE2294 || \
                   CYGPKG_HAL_ARM_LPC2XXX_OLPCH2294 || \
                   CYGPKG_HAL_ARM_LPC2XXX_OLPCL2294)

    requires      CYGPKG_DEVS_FLASH_STRATA_V2

    implements    CYGHWR_IO_FLASH_BLOCK_LOCKING

    description "
        Olimex LPC-X2294 boards all have strata family 28FxxxC3 flash
        memory parts. These parts have boot blocks. There is no buffered
        write capability. Individual blocks can be locked and unlocked
        in software"

}

