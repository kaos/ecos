# ====================================================================
#
#      hal_i386_pcmb.cdl
#
#      PC Motherboard HAL package configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  jskov
# Contributors:   nickg
# Date:           1999-11-01
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_I386_PCMB {
    display  "i386 PC Motherboard Support"
    parent        CYGPKG_HAL_I386
    define_header hal_i386_pcmb.h
    include_dir   cyg/hal
    description   "
    The i386 PC Motherboard HAL package provides the
    support needed to run eCos binaries on an i386 PC
    using a standard motherboard. This package provides
    support for the standard PC devices: timers, interrupt
    controller, serial ports, ASCII display, keyboard, PCI
    bus etc. that are found on all PC compatible platforms.
    It does not provide support for devices that may also be
    found on modern motherboards, such as ethernet, sound and
    video devices. These are supported by drivers elsewhere."

    compile      pcmb_misc.c pcmb_serial.c 

    implements   CYGINT_HAL_I386_MEM_REAL_REGION_TOP
    implements   CYGINT_HAL_PLF_IF_IDE
    
    # Real-time clock/counter specifics
    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants."
        description   "The RTC period is based on the clock input
	               to the 8254, which is 1193180 Hz.
	               CYGNUM_HAL_RTC_PERIOD is set for 100 ticks
	               per second."
        flavor        none
    
        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            calculated    1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            calculated    100
        }
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
           calculated     11932
        }
    }

    cdl_component CYGPKG_HAL_I386_PCMB_MEMSIZE {
        display       "How to discover the size of available RAM."
        flavor        data
        legal_values  {"BIOS" "HARDCODE"}
        default_value {"BIOS"}
        description   "It is possible for the HAL to discover the 
                       size of RAM In several ways. Currently this
                        can be done by querying the BIOS or by 
                        hardcoding the values into the executable."
 
        cdl_option CYGNUM_HAL_I386_PCMB_MEMSIZE_BASE {
            display       "Amount of Base RAM available."
            flavor        data
            default_value 0x000F0000
            active_if     { CYGPKG_HAL_I386_PCMB_MEMSIZE == "HARDCODE" }
        }
 
        cdl_option CYGNUM_HAL_I386_PCMB_MEMSIZE_EXTENDED {
            display       "Amount of Extended RAM available."
            flavor        data
            default_value 0x00100000
            active_if     { CYGPKG_HAL_I386_PCMB_MEMSIZE == "HARDCODE" }
        }
    }
 
    
    cdl_interface CYGINT_HAL_I386_PCMB_SCREEN_SUPPORT {
	display       "Enable PC screen support"
	compile       pcmb_screen.c
	description   "This option enables support for the PC screen and
	               keyboard. These are combined into a virtual serial
	               device that may be used for diagnostic output.
	               Note that there is little point in trying to use it
	               as a debug channel."
    }
}
