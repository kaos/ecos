#==========================================================================
# 
#       kbd_ipaq.cdl
# 
#       eCos configuration data for the Compaq iPAQ keypad/buttons
# 
#==========================================================================
#####COPYRIGHTBEGIN####
#                                                                           
#  The contents of this file are subject to the Red Hat eCos Public License 
#  Version 1.1 (the "License"); you may not use this file except in         
#  compliance with the License.  You may obtain a copy of the License at    
#  http://www.redhat.com/                                                   
#                                                                           
#  Software distributed under the License is distributed on an "AS IS"      
#  basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
#  License for the specific language governing rights and limitations under 
#  the License.                                                             
#                                                                           
#  The Original Code is eCos - Embedded Configurable Operating System,      
#  released September 30, 1998.                                             
#                                                                          
#  The Initial Developer of the Original Code is Red Hat.                   
#  Portions created by Red Hat are                                          
#  Copyright (C) 2001 Red Hat, Inc.
#  All Rights Reserved.                                                     
#                                                                           
#####COPYRIGHTEND####
#==========================================================================
######DESCRIPTIONBEGIN####
# 
# Author(s):    gthomas
# Contributors: gthomas
# Date:         2001-03-15
# Purpose:      
# Description:  Kbdscreen drivers for Compaq iPAQ
# 
#####DESCRIPTIONEND####
# 
#==========================================================================

cdl_package CYGPKG_DEVS_KBD_IPAQ {
    display     "Keypad driver for iPAQ"
    include_dir cyg/io

    active_if   CYGPKG_IO_FILEIO
    requires    CYGPKG_IO
    requires    CYGFUN_KERNEL_API_C
    requires    CYGPKG_HAL_ARM_SA11X0_IPAQ
    active_if   !CYGSEM_IPAQ_LCD_COMM

    compile       -library=libextras.a ipaq_kbd.c

    description "Keypad driver for the iPAQ using the Atmel micro-controller"

    cdl_component CYGPKG_DEVS_KBD_IPAQ_OPTIONS {
        display "options"
        flavor  none
        no_define

        cdl_option CYGPKG_DEVS_KBD_IPAQ_CFLAGS {
            display       "Additional compiler flags"
            flavor        data
            no_define
            default_value { "" }
            description "
               This option modifies the set of compiler flags for
               building the keypad driver package. These flags
               are used in addition to the set of global flags."
        }

        cdl_option CYGDAT_DEVS_KBD_IPAQ_NAME {
            display "Device name for the keypad driver"
            flavor data
            default_value {"\"/dev/kbd\""}
            description " This option specifies the name of the keypad device"
        }

        cdl_option CYGNUM_DEVS_KBD_IPAQ_EVENT_BUFFER_SIZE {
            display "Number of events the driver can buffer"
            flavor data
            default_value { 32 }
            description "
                This option defines the size of the keypad device internal
            buffer. The cyg_io_read() function will return as many of these
            as there is space for in the buffer passed."
        }
    }
}
