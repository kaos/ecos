# ====================================================================
#
#      hal_mips_sim.cdl
#
#      MIPS SIM HAL package configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  bartv
# Contributors:
# Date:           1999-11-02
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_MIPS_SIM {
    display  "Minimal simulator"
    parent        CYGPKG_HAL_MIPS
    define_header hal_mips_sim.h
    include_dir   cyg/hal
    description   "
           The minimal simulator HAL package is provided for when only
           a simple simulation of the processor architecture is
           desired, as opposed to detailed simulation of any specific
           board. To use this minimal simulator the command
           `target sim --board=jmr3904pal' should be used from inside
           gdb. It is not possible to use any of the eCos device
           drivers when the simulator is running in this mode"

    compile       hal_diag.c platform.S plf_misc.c

    implements CYGINT_HAL_DEBUG_GDB_CTRLC_UNSUPPORTED

    cdl_option CYGBLD_HAL_TARGET_H {
        display "architecture header file"
        flavor data
        no_define
	define -file system.h CYGBLD_HAL_TARGET_H
        calculated { CYGPKG_HAL_MIPS_TX39 ? "<pkgconf/hal_mips_tx39.h>" :
                                            "<pkgconf/hal_mips_vr4300.h>"}
    }

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_mips_sim.h>"
    }

    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        legal_values  {"RAM"}
        default_value {"RAM"}
	no_define
	define -file system.h CYG_HAL_STARTUP
        description   "
            Only supports RAM startup."
    }

    # Real-time clock/counter specifics
    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants."
        flavor        none
    
        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            calculated    1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            calculated    100
        }
        # Isn't a nice way to handle freq requirement!
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
            calculated    999
        }
    }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        parent  CYGPKG_NONE
        description   "
	    Global build options including control over
	    compiler flags, linker flags and choice of toolchain."


        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { CYGPKG_HAL_MIPS_TX39 ? "mips-tx39-elf" : \
						   "mips64vr4300-elf" }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { CYGPKG_HAL_MIPS_TX39 ? "-Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority" : "-mgp32 -EB -Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority" }
            description   "
                This option controls the global compiler flags which
                are used to compile all packages by
                default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { CYGPKG_HAL_MIPS_TX39 ? "-g -nostdlib -Wl,--gc-sections -Wl,-static" : "-mgp32 -EB -g -nostdlib -Wl,--gc-sections -Wl,-static" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { CYGPKG_HAL_MIPS_TX39 ? "mips_tx39_sim_ram" :
                                            "mips_vr4300_sim_ram" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { CYGPKG_HAL_MIPS_TX39 ? "<pkgconf/mlt_mips_tx39_sim_ram.ldi>" :
                                                "<pkgconf/mlt_mips_vr4300_sim_ram.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { CYGPKG_HAL_MIPS_TX39 ? "<pkgconf/mlt_mips_tx39_sim_ram.h>" : 
                                                "<pkgconf/mlt_mips_vr4300_sim_ram.h>" }
        }
    }
}
