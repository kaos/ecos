# ====================================================================
#
#      interrupts.cdl
#
#      configuration data related to kernel interrupt handling
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      bartv
# Original data:  nickg
# Contributors:
# Date:           1999-06-13
#
#####DESCRIPTIONEND####
#
# ====================================================================

# NOTE: the choice of list vs table should not be two separate
# options. There is a single option which must have one of
# two legal values.
cdl_component CYGIMP_KERNEL_INTERRUPTS_DSRS {
    display       "Use delayed service routines (DSRs)"
    default_value 1
    description   "
        In eCos the recommended way to handle device interrupts is to
        do a minimum amount of work inside the low level interrupt
        handler itself, and instead do as much as possible in a
        Delayed Service Routine or DSR. If an application does not
        make use of DSRs directly or indirectly then it is possible
        to disable the DSR support completely, which reduces the
        overheads of context switches and interrupt handling. Note
        that the kernel real-time clock makes use of DSRs, as do many
        of the device drivers. "

    cdl_interface CYGINT_KERNEL_INTERRUPTS_DSRS {
        requires 1 == CYGINT_KERNEL_INTERRUPTS_DSRS
        no_define
    }

    # NOTE: the choice of list vs table should not be two separate
    # options. There is a single option which must have one of
    # two legal values.
    cdl_option CYGIMP_KERNEL_INTERRUPTS_DSRS_LIST {
        display       "Use linked lists for DSRs"
        default_value 1
        implements    CYGINT_KERNEL_INTERRUPTS_DSRS
        description   "
            When DSR support is enabled the kernel must keep track of all
            the DSRs that are pending. This information can be kept in a
            fixed-size table or in a linked list. The list implementation
            requires that the kernel disable interrupts for a very short
            period of time outside interrupt handlers, but there is no
            possibility of a table overflow occurring."
    }

    cdl_component CYGIMP_KERNEL_INTERRUPTS_DSRS_TABLE {
        display       "Use fixed-size table for DSRs"
        default_value 0
        implements    CYGINT_KERNEL_INTERRUPTS_DSRS
        description   "
            When DSR support is enabled the kernel must keep track of all
            the DSRs that are pending. This information can be kept in a
            fixed-size table or in a linked list. The table
            implementation involves a very small risk of overflow at
            run-time if a given interrupt source is able to have more
            than one pending DSR. However it has the advantage that
            the kernel does not need to disable interrupts outside
            interrupt handlers."

        cdl_option CYGNUM_KERNEL_INTERRUPTS_DSRS_TABLE_SIZE {
            display       "Number of entries in fixed-size DSR table"
            flavor        data
            legal_values  2 to 1024
            default_value 32
            description "
            When DSR support is enabled the kernel must keep track of all
            the DSRs that are pending. One approach involves a fixed-size
            table, which involves a very small risk of overflow at
            run-time. By increasing the table size it is possible to reduce
            this risk."
        }
    }

    cdl_option CYGIMP_KERNEL_INTERRUPTS_CHAIN {
        display       "Chain all interrupts together"
        requires      CYGIMP_HAL_COMMON_INTERRUPTS_CHAIN
        default_value 0
        description "
            Interrupts can be attached to vectors either singly, or be
            chained together. The latter is necessary if there is no way
            of discovering which device has interrupted without
            inspecting the device itself. It can also reduce the amount
            of RAM needed for interrupt decoding tables and code."
    }
}
