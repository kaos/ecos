# ====================================================================
#
#      debugging.cdl
#
#      HAL debugging configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  nickg,jskov,jlarmour
# Contributors:
# Date:           1999-07-02
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_interface CYGINT_HAL_DEBUG_GDB_STUBS {
    display       "Support for GDB stubs"
    no_define
    description   "
        The HAL implements GDB stubs for the target."
}

cdl_option CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS {
    display       "Include GDB stubs in HAL"
    active_if     CYGINT_HAL_DEBUG_GDB_STUBS
    default_value 0
    requires      ! CYGSEM_HAL_USE_ROM_MONITOR
    description   "
        This option causes a set of GDB stubs to be included into the
        system. On some target systems the GDB support will be
        provided by other means, for example by a ROM monitor. On
        other targets, especially when building a ROM-booting system,
        the necessary support has to go into the target library
        itself."
}

cdl_interface CYGINT_HAL_DEBUG_GDB_STUBS_BREAK {
    display       "Support for external break support in GDB stubs"
    no_define
    description   "
        The HAL implements external break (or asynchronous interrupt)
        in the GDB stubs for the target."  
}

cdl_option CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT {
    display       "Include GDB external break support for stubs"
    active_if     CYGINT_HAL_DEBUG_GDB_STUBS_BREAK
    requires      CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
    default_value 0
    description   "
        This option causes the GDB stub to add a serial interrupt handler
        which will listen for GDB break packets. This lets you stop the
        target asynchronously when using GDB, usually by hitting Control+C
        or pressing the STOP button. This option differs from
        CYGDBG_HAL_DEBUG_GDB_CTRLC_SUPPORT in that it is used when
        GDB stubs are present."
}

cdl_interface CYGINT_HAL_DEBUG_GDB_CTRLC_UNSUPPORTED {
    display "Platform does not support CTRLC"
    no_define
}

cdl_option CYGDBG_HAL_DEBUG_GDB_CTRLC_SUPPORT {
    display       "Include GDB external break support when no stubs"
    requires      !CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT
    active_if     { CYGINT_HAL_DEBUG_GDB_CTRLC_UNSUPPORTED == 0 }
    default_value 1
    description   "
        This option adds an interrupt handler for the GDB serial line
        which will listen for GDB break packets. This lets you stop the
        target asynchronously when using GDB, usually by hitting Control+C
        or pressing the STOP button. This option differs from
        CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT in that it is used when the GDB
        stubs are NOT present."
}

cdl_option CYGDBG_HAL_DEBUG_GDB_THREAD_SUPPORT {
    display       "Include GDB multi-threading debug support"
    active_if     { CYGSEM_HAL_ROM_MONITOR || CYGDBG_KERNEL_DEBUG_GDB_THREAD_SUPPORT }
    default_value 1
    description   "
        This option enables some extra HAL code which is needed
        to support multi-threaded source level debugging."

    compile dbg-threads-syscall.c
}
