# ====================================================================
#
#      hal_arm_at91_eb42.cdl
#
#      ARM AT91 EB42 HAL package configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
## Copyright (C) 2003 Nick Garnett <nickg@calivar.com>
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Contributors:   gthomas, tkoeller, tdrury, nickg
# Date:           2001-07-12
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_ARM_AT91_EB42 {
    display       "Atmel EB42 eval board HAL"
    parent        CYGPKG_HAL_ARM_AT91
    define_header hal_arm_at91_eb42.h
    include_dir   cyg/hal
    hardware
    description   "
        The EB42 HAL package provides the support needed to run
        eCos on an Atmel EB42 eval board."

    compile       eb42_misc.c

    requires      { CYGHWR_HAL_ARM_AT91 == "M42800A" }

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H   <pkgconf/hal_arm.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_VARIANT_H  <pkgconf/hal_arm_at91.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_arm_at91_eb42.h>"
	puts $::cdl_header "#define HAL_PLATFORM_CPU    \"ARM7TDMI\""
        puts $::cdl_header "#define HAL_PLATFORM_BOARD  \"Atmel AT91/EB42\""
        puts $::cdl_header "#define HAL_PLATFORM_EXTRA  \"\""
    }

    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        default_value {"RAM"}
        legal_values  {"RAM" "ROM" "ROMRAM"}
	no_define
	define -file system.h CYG_HAL_STARTUP
        description   "
            When targetting the EB42 eval board it is possible to build
            the system for either RAM bootstrap or ROM bootstrap(s). Select
            'ram' when building programs to load into RAM using onboard
            debug software such as Angel or eCos GDB stubs.  Select 'rom'
            when building a stand-alone application which will be put
            into ROM.  Using ROMRAM will allow the program to exist in
            ROM, but be copied to RAM during startup."
    }

    # Real-time clock/counter specifics
    cdl_option CYGNUM_HAL_ARM_AT91_CLOCK_SPEED {
        display       "CPU clock speed"
        flavor        data
        calculated    32768000
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
        display      "Number of communication channels on the board"
        flavor       data
        calculated   2
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
        display          "Debug serial port"
        active_if        CYGPRI_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_CONFIGURABLE
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
            The EB42 board has two serial ports. This option
            chooses which port will be used to connect to a host
            running GDB."
     }

     cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
         display          "Diagnostic serial port"
         active_if        CYGPRI_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_CONFIGURABLE
         flavor data
         legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
         default_value    0
         description      "
            The EB42 board has two serial ports. This option
            chooses which port will be used for diagnostic output."
     }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CHANNELS_DEFAULT_BAUD {
        display       "Console/GDB serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 57600 115200
        default_value 38400
        description   "
            This option controls the default baud rate used for the
            Console/GDB connection."
    }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        parent  CYGPKG_NONE
        description   "
	    Global build options including control over
	    compiler flags, linker flags and choice of toolchain."


        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "arm-elf" }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { "-mcpu=arm7tdmi -mno-short-load-words -Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority" }
            description   "
                This option controls the global compiler flags which are used to
                compile all packages by default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { "-mcpu=arm7tdmi -mno-short-load-words -Wl,--gc-sections -Wl,-static -g -nostdlib" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { (CYG_HAL_STARTUP == "RAM") ?    "arm_at91_eb42_ram" :
                     (CYG_HAL_STARTUP == "ROMRAM") ? "arm_at91_eb42_romram" :
                                                     "arm_at91_eb42_rom" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { (CYG_HAL_STARTUP == "RAM") ? "<pkgconf/mlt_arm_at91_eb42_ram.ldi>" :
                         (CYG_HAL_STARTUP == "ROMRAM") ? "<pkgconf/mlt_arm_at91_eb42_romram.ldi>" :
                                                      "<pkgconf/mlt_arm_at91_eb42_rom.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { (CYG_HAL_STARTUP == "RAM") ? "<pkgconf/mlt_arm_at91_eb42_ram.h>" :
                         (CYG_HAL_STARTUP == "ROMRAM") ? "<pkgconf/mlt_arm_at91_eb42_romram.h>" :
                                                      "<pkgconf/mlt_arm_at91_eb42_rom.h>" }
        }
    }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "ROM" || CYG_HAL_STARTUP == "ROMRAM" }
        description   "
            Enable this option if this program is to be used as a ROM monitor,
            i.e. applications will be loaded into RAM on the board, and this
            ROM monitor may process exceptions or interrupts generated from the
            application. This enables features such as utilizing a separate
            interrupt stack when exceptions are generated."
    }

    cdl_option CYGSEM_HAL_USE_ROM_MONITOR {
         display       "Work with a ROM monitor"
         flavor        booldata
         legal_values  { "Generic" "GDB_stubs" }
         default_value { CYG_HAL_STARTUP == "RAM" ? "GDB_stubs" : 0 }
         parent        CYGPKG_HAL_ROM_MONITOR
         requires      { CYG_HAL_STARTUP == "RAM" }
         description   "
             Support can be enabled for different varieties of ROM monitor.
             This support changes various eCos semantics such as the encoding
             of diagnostic output, or the overriding of hardware interrupt
             vectors.
             Firstly there is \"Generic\" support which prevents the HAL
             from overriding the hardware vectors that it does not use, to
             instead allow an installed ROM monitor to handle them. This is
             the most basic support which is likely to be common to most
             implementations of ROM monitor.
             \"GDB_stubs\" provides support when GDB stubs are included in
             the ROM monitor or boot ROM."
     }

    cdl_component CYGPKG_REDBOOT_HAL_OPTIONS {
        display       "Redboot HAL options"
        flavor        none
        no_define
        parent        CYGPKG_REDBOOT
        active_if     CYGPKG_REDBOOT
        description   "
            This option lists the target's requirements for a valid Redboot
            configuration."

        cdl_option CYGBLD_BUILD_REDBOOT_BIN {
            display       "Build Redboot ROM binary image"
            active_if     CYGBLD_BUILD_REDBOOT
            default_value 1
            no_define
            description "This option enables the conversion of the Redboot ELF
                         image to a binary image suitable for ROM programming."

            make -priority 325 {
                <PREFIX>/bin/redboot.bin : <PREFIX>/bin/redboot.elf
                $(OBJCOPY) --strip-debug $< $(@:.bin=.img)
                $(OBJCOPY) -O srec $< $(@:.bin=.srec)
                $(OBJCOPY) -O binary $< $@
            }

        }
    }
}
