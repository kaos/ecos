# ====================================================================
#
#      ser_mips_jmr3904.cdl
#
#      eCos serial MIPS/JMR3904 configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  gthomas
# Contributors:
# Date:           1999-07-14
#
#####DESCRIPTIONEND####
#
# ====================================================================


cdl_package CYGPKG_IO_SERIAL_TX39_JMR3904 {
    display       "TX39 JMR3904 serial device drivers"

    parent        CYGPKG_IO_SERIAL_DEVICES
    active_if     CYGPKG_IO_SERIAL
    active_if     CYGPKG_HAL_MIPS_TX39_JMR3904

    requires      CYGPKG_ERROR
    include_dir   cyg/io
#    include_files ; # none _exported_ whatsoever
    description   "
           This option enables the serial device drivers for the
           TX39 JMR3904."
    doc           redirect/ecos-device-drivers.html

    compile       -library=libextras.a   tx3904_serial.c

    define_proc {
        puts $::cdl_system_header "/***** serial driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_DEVICE_HEADER <pkgconf/io_serial_tx39_jmr3904.h>"
        puts $::cdl_system_header "/*****  serial driver proc output end  *****/"
    }

# FIXME: Bad name
cdl_option CYGPKG_IO_SERIAL_TX39_JMR3904_POLLED_MODE {
    display       "TX39 JMR3904 polled mode serial drivers"
    flavor        bool
    default_value 0
    description   "
        If asserted, this option specifies that the serial device
        drivers for the TX39 JMR3904 should be polled-mode instead of
        interrupt driven."
}

cdl_component CYGPKG_IO_SERIAL_TX39_JMR3904_SERIAL0 {
    display       "TX39 JMR3904 serial port 0 driver"
    flavor        bool
    default_value 1
    description   "
        This option includes the serial device driver for port 0 on the 
        TX39 JMR3904."

    cdl_option CYGDAT_IO_SERIAL_TX39_JMR3904_SERIAL0_NAME {
        display       "Device name for TX39 JMR3904 serial port 0"
        flavor        data
        default_value {"\"/dev/ser0\""}
        description   "
            This option specifies the device name port 0 on the TX39 JMR3904."
    }

    cdl_option CYGNUM_IO_SERIAL_TX39_JMR3904_SERIAL0_BAUD {
        display       "Baud rate for the TX39 JMR3904 serial port 0 driver"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 234000
        }
        default_value 38400
        description   "
            This option specifies the default baud rate (speed) for the 
            TX39 JMR3904 port 0."
    }

    cdl_option CYGNUM_IO_SERIAL_TX39_JMR3904_SERIAL0_BUFSIZE {
        display       "Buffer size for the TX39 JMR3904 serial port 0 driver"
        flavor        data
        legal_values  0 to 8192
        default_value 128
        description   "
            This option specifies the size of the internal buffers used
            for the TX39 JMR3904 port 0."
    }
}
cdl_component CYGPKG_IO_SERIAL_TX39_JMR3904_SERIAL1 {
    display       "TX39 JMR3904 serial port 1 driver"
    flavor        bool
    default_value 1
    description   "
        This option includes the serial device driver for port 1 on 
        the TX39 JMR3904."

    cdl_option CYGDAT_IO_SERIAL_TX39_JMR3904_SERIAL1_NAME {
        display       "Device name for TX39 JMR3904 serial port 1"
        flavor        data
        default_value {"\"/dev/ser1\""}
        description   "
            This option specifies the device name port 1 on the TX39 JMR3904."
    }

    cdl_option CYGNUM_IO_SERIAL_TX39_JMR3904_SERIAL1_BAUD {
        display       "Baud rate for the TX39 JMR3904 serial port 1 driver"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 234000
        }
        default_value 38400
        description   "
            This option specifies the default baud rate (speed) for the
            TX39 JMR3904 port 1."
    }

    cdl_option CYGNUM_IO_SERIAL_TX39_JMR3904_SERIAL1_BUFSIZE {
        display       "Buffer size for the TX39 JMR3904 serial port 1 driver"
        flavor        data
        legal_values  0 to 8192
        default_value 128
        description   "
            This option specifies the size of the internal buffers used 
            for the TX39 JMR3904 port 1."
    }
}

    cdl_component CYGPKG_IO_SERIAL_MIPS_JMR3904_OPTIONS {
        display "Serial device driver build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_IO_SERIAL_MIPS_JMR3904_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_IO_SERIAL_MIPS_JMR3904_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are removed from
                the set of global flags if present."
        }
    }
}

# EOF ser_mips_jmr3904.cdl
