# ====================================================================
#
#      hal_powerpc_ppc60x.cdl
#
#      PowerPC/PPC60x variant architectural HAL package configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Contributors:
# Date:           2000-02-04
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_POWERPC_PPC60x {
    display       "PowerPC 60x variant HAL"
    parent        CYGPKG_HAL_POWERPC
    hardware
    include_dir   cyg/hal
    define_header hal_powerpc_ppc60x.h
    description   "
           The PowerPC 60x variant HAL package provides generic support
           for this processor variant. It is also necessary to
           select a specific target platform HAL package."

    # Note: This should be sub-variant specific to reduce memory use.
    define_proc {
        puts $cdl_header "#define CYGHWR_HAL_VSR_TABLE (CYGHWR_HAL_POWERPC_VECTOR_BASE + 0x3000)"
        puts $cdl_header "#define CYGHWR_HAL_VIRTUAL_VECTOR_TABLE (CYGHWR_HAL_VSR_TABLE + 0x200)"
    }

    cdl_component CYGPKG_HAL_POWERPC_PPC603 {
        display       "PowerPC 603 microprocessor"
        default_value 1
        implements    CYGINT_HAL_POWERPC_VARIANT
        description "
            The PowerPC 603 microprocessor."

        cdl_option CYGHWR_HAL_POWERPC_FPU {
            display    "Variant FPU support"
            calculated 1
        }

        cdl_option CYGPKG_HAL_POWERPC_MSBFIRST {
            display    "CPU Variant big-endian"
            calculated 1
        }
    }

    define_proc {
        puts $::cdl_header "#include <pkgconf/hal_powerpc.h>"
    }

    compile       var_intr.c var_misc.c variant.S
}
