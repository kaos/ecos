# ====================================================================
#
#      smsc_lan91cxx_eth_drivers.cdl
#
#      Ethernet drivers - support for LAN91CXX compatible ethernet controllers
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Contributors:   gthomas, jskov
# Date:           2000-11-22
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_SMSC_LAN91CXX {
    display       "SMSC LAN91CXX compatible ethernet driver"
    description   "Ethernet driver for SMSC LAN91CXX compatible controllers."

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_IO_ETH_DRIVERS

    active_if     CYGINT_DEVS_ETH_SMSC_LAN91CXX_REQUIRED

    include_dir   .
    include_files ; # none _exported_ whatsoever
    compile       -library=libextras.a if_lan91cxx.c

    define_proc {
        puts $::cdl_header "#include <pkgconf/system.h>";
        puts $::cdl_header "#include CYGDAT_DEVS_ETH_SMSC_LAN91CXX_CFG";
    }

    cdl_option CYGSEM_DEVS_ETH_SMSC_LAN91CXX_WRITE_EEPROM {
	display "SIOCSIFHWADDR records ESA (MAC address) in EEPROM"
	default_value 0
	description   "
	    The ioctl() socket call with operand SIOCSIFHWADDR sets the
	    interface hardware address - the MAC address or Ethernet Station
	    Address (ESA).  This option causes the new MAC address to be written
	    into the EEPROM associated with the interface, so that the new
	    MAC address is permanently recorded.  Doing this should be a
	    carefully chosen decision, hence this option."
    }

    cdl_interface CYGINT_DEVS_ETH_SMSC_LAN91CXX_STATIC_ESA {
	display "ESA is statically configured"
	description "
	    If this is nonzero, then the ESA (MAC address) is statically
            configured in the platform-specific package which instantiates
	    this driver with all its details."
    }

    cdl_interface CYGINT_DEVS_ETH_SMSC_LAN91CXX_PCMCIA_MODE {
	display "Chip is wired in PCMCIA mode"
	description "
	    If this is nonzero, then the chip is assumed to be hardware
            configured in PCMCIA mode."
    }

    cdl_component CYGPKG_DEVS_ETH_SMSC_LAN91CXX_OPTIONS {
        display "LAN91CXX ethernet driver build options"
        flavor  none
	no_define

        cdl_option CYGPKG_DEVS_ETH_SMSC_LAN91CXX_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building the LAN91CXX ethernet driver package.
                These flags are used in addition
                to the set of global flags."
        }
    }
}
