# ====================================================================
#
#      ser_sh_edk7708.cdl
#
#      eCos serial SH/EDK7708 configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Contributors:
# Date:           1999-07-08
#
#####DESCRIPTIONEND####
#
# ====================================================================


cdl_package CYGPKG_IO_SERIAL_SH_EDK7708 {
    display       "SH3 EDK7708  serial device drivers"

    parent        CYGPKG_IO_SERIAL_DEVICES
    active_if     CYGPKG_IO_SERIAL
    active_if     CYGPKG_HAL_SH_EDK7708

    requires      CYGPKG_ERROR
    include_dir   cyg/io
    include_files ; # none _exported_ whatsoever
    description   "
           This option enables the serial device drivers for the
           Hitachi SH3 EDK7708 board."
    doc           redirect/ecos-device-drivers.html


    define_proc {
        puts $::cdl_system_header "/***** serial driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_DEVICE_HEADER <pkgconf/io_serial_sh_edk7708.h>"
        puts $::cdl_system_header "/*****  serial driver proc output end  *****/"
    }

cdl_component CYGPKG_IO_SERIAL_SH_EDK7708_SCI {
    display       "SH3 EDK7708 SCI device driver"
    flavor        bool
    default_value 1
    description   "
        This option includes the serial device driver for the SCI port."

    compile       -library=libextras.a   sh_sci_serial.c

    cdl_option CYGDAT_IO_SERIAL_SH_EDK7708_SCI_NAME {
        display       "Device name for SH3 EDK7708 SCI"
        flavor        data
        default_value {"\"/dev/ser1\""}
        description   "
            This option specifies the device name for the SCI port."
    }

    cdl_option CYGNUM_IO_SERIAL_SH_EDK7708_SCI_BAUD {
        display       "Baud rate for the SH SCI driver"
        flavor        data
        legal_values  { 4800 9600 14400 19200 38400 57600 115200 }
        default_value 38400
        description   "
            This option specifies the default baud rate (speed) for the 
            SCI port."
    }

    cdl_option CYGNUM_IO_SERIAL_SH_EDK7708_SCI_BUFSIZE {
        display       "Buffer size for the SH SCI driver"
        flavor        data
        legal_values  0 to 8192
        default_value 128
        description   "
            This option specifies the size of the internal buffers used for
            the SCI port."
    }
}

    cdl_component CYGPKG_IO_SERIAL_SH_EDK7708_OPTIONS {
        display "Serial device driver build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_IO_SERIAL_SH_EDK7708_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_IO_SERIAL_SH_EDK7708_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are removed from
                the set of global flags if present."
        }
    }
}

# EOF ser_sh_edk7708.cdl
