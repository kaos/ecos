# ====================================================================
#
#      hal_mn10300_am33_asb2305.cdl
#
#      AM33-2/ASB2305 board HAL package configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
# -------------------------------------------
# This file is part of eCos, the Embedded Configurable Operating System.
# Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
#
# eCos is free software; you can redistribute it and/or modify it under
# the terms of the GNU General Public License as published by the Free
# Software Foundation; either version 2 or (at your option) any later version.
#
# eCos is distributed in the hope that it will be useful, but WITHOUT ANY
# WARRANTY; without even the implied warranty of MERCHANTABILITY or
# FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
# for more details.
#
# You should have received a copy of the GNU General Public License along
# with eCos; if not, write to the Free Software Foundation, Inc.,
# 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
#
# As a special exception, if other files instantiate templates or use macros
# or inline functions from this file, or you compile this file and link it
# with other works to produce a work based on this file, this file does not
# by itself cause the resulting work to be covered by the GNU General Public
# License. However the source code for this file must still be made available
# in accordance with section (3) of the GNU General Public License.
#
# This exception does not invalidate any other reasons why a work based on
# this file might be covered by the GNU General Public License.
#
# Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
# at http://sources.redhat.com/ecos/ecos-license
# -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      dhowells
# Original data:  dmoseley. nick, bartv
# Contributors:
# Date:           2001-05-17
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_MN10300_AM33_ASB2305 {
    display  "Panasonic ASB2305 Evaluation Board"
    parent        CYGPKG_HAL_MN10300
    requires      CYGPKG_HAL_MN10300_AM33
    requires      { CYGHWR_HAL_MN10300_AM33_REVISION == 2 }
    define_header hal_mn10300_am33_asb2305.h
    include_dir   cyg/hal
    description   "
           The ASB2305 HAL package should be used when targetting the
           actual hardware for the Panasonic ASB2305 Evaluation Board
           with the MN103E010 microcontroller."

    compile       hal_diag.c plf_stub.c plf_misc.c ser_asb.c

    implements    CYGINT_HAL_DEBUG_GDB_STUBS
    implements    CYGINT_HAL_DEBUG_GDB_STUBS_BREAK
    implements    CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT

    requires CYGSEM_HAL_UNCACHED_FLASH_ACCESS == 1;

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H   <pkgconf/hal_mn10300_am33.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_mn10300_am33_asb2305.h>"
        puts $::cdl_system_header "#define HAL_PLATFORM_BOARD    \"Panasonic ASB2305\""
        puts $::cdl_system_header "#define HAL_PLATFORM_EXTRA    \"\""
        puts $::cdl_system_header "#define HAL_PLATFORM_CPU      \"MN103E010 AM33/2.0\""
    }

    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        legal_values  {"RAM" "ROM"}
        default_value {"ROM"}
        no_define
        define -file system.h CYG_HAL_STARTUP
        description   "
            This determines whether the stored .data section will need copying
            to RAM before it can be used."
    }

    cdl_component CYG_HAL_ROM_SLOT {
        display       "ROM slot in which residing"
        flavor        data
        legal_values  {"BootPROM" "SysFlash"}
        default_value {"BootPROM"}
        no_define
        define -file system.h CYG_HAL_ROM_SLOT
        description   "
            This specifies which ROM slot the program resides in (and is booted
            from."
    }

    # Real-time clock/counter specifics
    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants."
        description   "
            The NUMERATOR divided by the DENOMINATOR gives the number of
            nanoseconds per tick. The PERIOD is the divider to be programmed
            into a hardware timer that is driven from an appropriate hardware
            clock, such that the timer overflows once per tick (normally
            generating a CPU interrupt to mark the end of a tick). The tick
            rate is typically 100Hz.
            The clock is generated with onboard 16-bit timers TM4 and TM5
            cascaded together to form a 32-bit timer."
        flavor none

        cdl_option CYGHWR_HAL_MN10300_IOCLK_SPEED {
            display          "Processor I/O clock speed (Hz)"
            flavor           data
            calculated       (25 * 1000 * 1000)
            description      "
                The processor I/O clock speed, from which onboard timers can
                draw their sources."
        }

        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            calculated    (1000 * 1000 * 1000)
        }

        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            calculated    100
        }

        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock divisor"
            flavor        data
            calculated    (CYGHWR_HAL_MN10300_IOCLK_SPEED * CYGNUM_HAL_RTC_NUMERATOR) / (1000000000 * CYGNUM_HAL_RTC_DENOMINATOR)
        }
    }

    cdl_option CYGHWR_HAL_MN10300_AM33_ASB_DIAG_PORT {
        display          "Diagnostic Serial Port"
        flavor data
        legal_values     0 1
        default_value    0
        description      "
           The ASB2305 board has two serial ports. This option
           chooses which of these ports will be used for diagnostic output.
           At present only port 0 is supported."
   }

   cdl_option CYGHWR_HAL_MN10300_AM33_ASB_DIAG_BAUD {
       display          "Diagnostic Serial Port Baud Rate"
       flavor data
       legal_values     9600 19200 38400 115200
       default_value    38400
       description      "
           This option selects the baud rate used for the diagnostic port.
           Note: this should match the value chosen for the GDB port if the
           diagnostic and GDB port are the same."
   }

   cdl_option CYGHWR_HAL_MN10300_AM33_ASB_GDB_PORT {
       display          "GDB Serial Port"
       flavor data
       legal_values     0 1
       default_value    0
       description      "
           The ASB2305 board has two separate serial ports.  This option
           chooses which of these ports will be used to connect to a host
           running GDB.
           At present only port 0 is supported."
   }

   cdl_option CYGHWR_HAL_MN10300_AM33_ASB_GDB_BAUD {
       display          "GDB Serial Port Baud Rate"
       flavor data
       legal_values     9600 19200 38400 115200
       default_value    38400
       description      "
           This option controls the baud rate used for the GDB connection."
   }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        parent  CYGPKG_NONE
        description   "
            Global build options including control over
            compiler flags, linker flags and choice of toolchain."


        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "mn10300-elf" }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { "-mam33-2 -Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -Wp,-Wno-paste -g -O2 -fno-builtin -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority" }
            description   "
                This option controls the global compiler flags which
                are used to compile all packages by
                default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { "-mam33 -g -nostdlib -Wl,--gc-sections -Wl,-static" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }

        cdl_option CYGBLD_BUILD_GDB_STUBS {
            display "Build GDB stub ROM image"
            default_value 0
            requires { CYG_HAL_STARTUP == "ROM" }
            requires CYGSEM_HAL_ROM_MONITOR
            requires CYGBLD_BUILD_COMMON_GDB_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
            requires ! CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT
            requires ! CYGDBG_HAL_DEBUG_GDB_THREAD_SUPPORT
            requires ! CYGDBG_HAL_COMMON_INTERRUPTS_SAVE_MINIMUM_CONTEXT
            requires ! CYGDBG_HAL_COMMON_CONTEXT_SAVE_MINIMUM
            no_define
            description "
                This option enables the building of the GDB stubs for the
                board. The common HAL controls takes care of most of the
                build process, but the final conversion from ELF image to
                binary data is handled by the platform CDL, allowing
                relocation of the data if necessary."

            make -priority 320 {
                <PREFIX>/bin/gdb_module.bin : <PREFIX>/bin/gdb_module.img
                $(OBJCOPY) -O binary $< $@
            }
        }
    }

    cdl_option CYGNUM_HAL_BREAKPOINT_LIST_SIZE {
        display       "Number of breakpoints supported by the HAL."
        flavor        data
        default_value 25
        description   "
            This option determines the number of breakpoints supported by the HAL."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
        display      "Number of communication channels on the board"
        flavor       data
        calculated   1
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
        display          "Debug serial port"
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
           The ASB2305 board has two serial ports.  Currently,
           only the first serial port is supported. This option
           chooses which port will be used to connect to a host
           running GDB."
    }

     cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
        display          "Diagnostic serial port"
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
           The ASB2305 board has two serial ports. Currently,
           only the first serial port is supported. This option
           chooses which port will be used for diagnostic output."
     }

     cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD {
        display          "Diagnostic serial port baudrates"
        flavor data
        legal_values     9600 19200 38400 57600 115200
        default_value    38400
        description      "
           The ASB2305 debug serial port baud rate setting."
     }

     cdl_option CYGSEM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_RTSCTS {
        display          "Diagnostic serial port RTS/CTS flow control"
        flavor           bool
        default_value    0
        description      "
           The ASB2305 debug serial port RTS/CTS flow control setting."
     }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { CYG_HAL_STARTUP  == "RAM"      ? "mn10300_am33_asb2305_ram" : \
                     CYG_HAL_ROM_SLOT == "BootPROM" ? "mn10300_am33_asb2305_rom" : \
                                                      "mn10300_am33_asb2305_flash" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { CYG_HAL_STARTUP == "RAM"       ? "<pkgconf/mlt_mn10300_am33_asb2305_ram.ldi>" : \
                         CYG_HAL_ROM_SLOT == "BootPROM" ? "<pkgconf/mlt_mn10300_am33_asb2305_rom.ldi>" : \
                                                          "<pkgconf/mlt_mn10300_am33_asb2305_flash.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { CYG_HAL_STARTUP == "RAM"       ? "<pkgconf/mlt_mn10300_am33_asb2305_ram.h>" : \
                         CYG_HAL_ROM_SLOT == "BootPROM" ? "<pkgconf/mlt_mn10300_am33_asb2305_rom.h>" : \
                                                          "<pkgconf/mlt_mn10300_am33_asb2305_flash.h>" }
        }
    }

    cdl_option CYGSEM_HAL_USE_ROM_MONITOR {
        display       "Work with a ROM monitor"
        flavor        booldata
        legal_values  { "GDB_stubs" }
        default_value { CYG_HAL_STARTUP == "RAM" ? "GDB_stubs" : 0 }
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "RAM" }
        description   "
            Support can be enabled for boot ROMs or ROM monitors which contain
            GDB stubs. This support changes various eCos semantics such as
            the encoding of diagnostic output, and the overriding of hardware
            interrupt vectors."
    }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 1
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "ROM" }
        description   "
            Enable this option if this program is to be used as a ROM monitor,
            i.e. applications will be loaded into RAM on the board, and this
            ROM monitor may process exceptions or interrupts generated from the
            application. This enables features such as utilizing a separate
            interrupt stack when exceptions are generated."
    }

    cdl_component CYGPKG_REDBOOT_HAL_OPTIONS {
        display       "Redboot HAL options"
        flavor        none
        no_define
        parent        CYGPKG_REDBOOT
        active_if     CYGPKG_REDBOOT
        description   "
            This option lists the target's requirements for a valid Redboot
            configuration."

        compile -library=libextras.a redboot_cmds.c

        cdl_option CYGBLD_BUILD_REDBOOT_BIN {
            display       "Build Redboot ROM binary image"
            active_if     CYGBLD_BUILD_REDBOOT
            default_value 1
            no_define
            description "This option enables the conversion of the Redboot ELF
                         image to a binary image suitable for ROM programming."
    
            make -priority 325 {
                <PREFIX>/bin/redboot.bin : <PREFIX>/bin/redboot.elf
                $(OBJCOPY) -O binary $< $@
            }
        }
    }
}
