# ====================================================================
#
#      hal_arm_xscale_verde.cdl
#
#      Intel XScale architectural HAL package configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      msalter
# Original data:  msalter
# Contributors:
# Date:           2001-12-03
#
#####DESCRIPTIONEND####
#
# ====================================================================
cdl_package CYGPKG_HAL_ARM_XSCALE_VERDE {
    display       "Intel XScale 80321 IO Processor"
    parent        CYGPKG_HAL_ARM
    hardware
    include_dir   cyg/hal
    define_header hal_arm_xscale_verde.h
    description   "
        This HAL variant package provides generic
        support for the Intel 80321 IO processors. It is also
        necessary to select a specific target platform HAL
        package."

    implements    CYGINT_HAL_ARM_ARCH_XSCALE

    # Let the architectural HAL see this variant's interrupts file
     define_proc {
        puts $::cdl_header \
       "#define CYGBLD_HAL_VAR_INTS_H <cyg/hal/hal_var_ints.h>"

        puts $::cdl_system_header "#define CYGBLD_HAL_ARM_VAR_IO_H"
    }

    compile       verde_misc.c verde_pci.c

    cdl_option CYGHWR_HAL_ARM_XSCALE_PROCESSOR_CCLK {
        display       "Processor clock rate"
        flavor        data
        default_value { CYGHWR_HAL_ARM_XSCALE_PROCESSOR_CCLK_DEFAULT ?
                        CYGHWR_HAL_ARM_XSCALE_PROCESSOR_CCLK_DEFAULT : 600000}
        description   "
           The XScale processor can run at various frequencies.
           These values are expressed in KHz."
    }

    # Real-time clock/counter specifics
    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants"
        flavor        none
        no_define
    
        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            calculated    1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            default_value 100
            description   "
              This option selects the heartbeat rate for the real-time clock.
              The rate is specified in ticks per second.  Change this value
              with caution - too high and your system will become saturated
              just handling clock interrupts, too low and some operations
              such as thread scheduling may become sluggish."
        }
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
            calculated    1000000/CYGNUM_HAL_RTC_DENOMINATOR
	    description   "
              This value gives the RTC period in microseconds. It is
              translated into the actual clock period value in the clock
              init and read functions."
        }
    }

    cdl_component CYGPKG_REDBOOT_XSCALE_OPTIONS {
        display       "Redboot for XScale options"
        flavor        none
        no_define
        parent        CYGPKG_REDBOOT
        active_if     CYGPKG_REDBOOT
        description   "
            This option lists the target's requirements for a valid Redboot
            configuration."

        # RedBoot details
        requires { CYGSEM_REDBOOT_ARM_LINUX_BOOT }
        requires { CYGHWR_REDBOOT_ARM_LINUX_EXEC_ADDRESS_DEFAULT == 0xc0008000 }
        define_proc {
            puts $::cdl_header "#define CYGHWR_REDBOOT_ARM_TRAMPOLINE_ADDRESS 0x00001f00"
        }
    }
}
