# ====================================================================
#
#      snmplib.cdl
#
#      SNMP library configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      hmt
# Original data:  hmt
# Contributors:   gthomas
# Date:           2000-05-30
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_SNMPLIB {
    display       "SNMP library"
    parent        CYGPKG_NET
#    doc           doc/index.html
    include_dir   ucd-snmp
    requires      CYGPKG_IO
    requires      { 0 != CYGINT_ISO_STRING_STRFUNCS }
    requires      { 0 != CYGINT_ISO_STRING_MEMFUNCS }
    requires      { 0 != CYGINT_ISO_STDLIB_STRCONV }
    requires      { 0 != CYGINT_ISO_STDIO_FORMATTED_IO }
    requires      { 0 != CYGINT_ISO_STRING_STRFUNCS }
    requires      { 0 != CYGINT_ISO_MALLOC }
    requires      { 0 != CYGINT_ISO_ERRNO }
    requires      { 0 != CYGINT_ISO_ERRNO_CODES }
    requires      CYGPKG_NET
    description   "SNMP protocol support library based on the UCD-SNMP project."

    compile					\
		asn1.c				\
		callback.c			\
		default_store.c			\
		int64.c				\
		keytools.c			\
		lcd_time.c			\
		md5.c				\
		mib.c				\
		mt_support.c			\
		parse.c				\
		read_config.c			\
		scapi.c				\
		snmp.c				\
		snmp_alarm.c			\
		snmp_api.c			\
		snmp_auth.c			\
		snmp_client.c			\
		snmp_debug.c			\
		snmp_logging.c			\
		snmpusm.c			\
		snmpv3.c			\
		system.c			\
		tools.c				\
		vacm.c


    cdl_option CYGDBG_NET_SNMPLIB_DEBUG {
	display        "Enable SNMP debug printout"
	flavor         bool
	default_value  0
	description "
	    This option enables the debugging printout facilities of the
	    UCD SNMP module, controlled by the global variable 'dodebug'.
	    Setting this variable produces lots of printout for SNMP agent
	    activity, often enough to make your SNMP client time out."
    }

    cdl_component CYGPKG_SNMPLIB_OPTIONS {
        display "SNMP library build options"
        flavor  none
	no_define

        cdl_option CYGPKG_SNMPLIB_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS -I$(PREFIX)/include/ucd-snmp" }
            description   "
                This option modifies the set of compiler flags for
                building the SNMP library package.
	        These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_SNMPLIB_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the SNMP library package. These flags are removed from
                the set of global flags if present."
        }
    }
}

# EOF snmplib.cdl
