# ====================================================================
#
#      startup.cdl
#
#      Infrastructure startup configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      bartv
# Original data:  bartv,hmt
# Contributors:
# Date:           1999-06-13
#
#####DESCRIPTIONEND####
#
# ====================================================================

# =================================================================
# The following options allow particular compatibility modes to be
# enabled, when they require specialised support from the startup
# process. These can affect the environment in which the program
# runs.
#
# CYGSEM_START_ISO_C_COMPATIBILITY enables compatibility with ISO C,
# in particular in eCos it creates a thread that invokes the function
# main() which the user must supply. It does this by invoking the function
# cyg_iso_c_start(). For more information, refer to the C library
# documentation.
#
# CYGSEM_START_UITRON_COMPATIBILITY enables compatibility with uItron.
# You must configure uItron with the correct tasks, and then enabling this
# option starts the uItron subsystem. It does this by invoking the function
# cyg_uitron_start().
#
# Both these can also be done by the user overriding cyg_user_start(),
# cyg_package_start(), or cyg_prestart(). Refer to the documentation on
# how and when to do this.

cdl_option CYGSEM_START_ISO_C_COMPATIBILITY {
    display       "Start ISO C library"
    default_value 1
    requires      CYGPKG_LIBC
    active_if     CYGPKG_LIBC
    description   "
        Generate a call to initialize the ISO C library
        (libc) within the system version of cyg_package_start().
        This enables compatibility with ISO C, in particular in
        eCos it creates a thread that invokes the function main()
        which the user must supply.
        It does this by invoking the function cyg_iso_c_start().
        If this is disabled, and you want to use the C library, you
        call cyg_iso_c_start() from your own cyg_package_start()
        or cyg_userstart()."
}
cdl_option CYGSEM_START_UITRON_COMPATIBILITY {
    display       "Start uITRON subsystem"
    default_value 0
    requires      CYGPKG_UITRON
    active_if     CYGPKG_UITRON
    description   "
        Generate a call to initialize the
        uITRON compatibility subsystem
        within the system version of cyg_package_start().
        This enables compatibility with uITRON.
        You must configure uITRON with the correct tasks before
        starting the uItron subsystem.
        If this is disabled, and you want to use uITRON,
        you must call cyg_uitron_start() from your own
        cyg_package_start() or cyg_userstart()."
}
