# ====================================================================
#
#      amd_pcnet_eth_drivers.cdl
#
#      Ethernet drivers - support for AMD PCNET ethernet controllers
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
# -------------------------------------------
# This file is part of eCos, the Embedded Configurable Operating System.
# Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
#
# eCos is free software; you can redistribute it and/or modify it under
# the terms of the GNU General Public License as published by the Free
# Software Foundation; either version 2 or (at your option) any later version.
#
# eCos is distributed in the hope that it will be useful, but WITHOUT ANY
# WARRANTY; without even the implied warranty of MERCHANTABILITY or
# FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
# for more details.
#
# You should have received a copy of the GNU General Public License along
# with eCos; if not, write to the Free Software Foundation, Inc.,
# 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
#
# As a special exception, if other files instantiate templates or use macros
# or inline functions from this file, or you compile this file and link it
# with other works to produce a work based on this file, this file does not
# by itself cause the resulting work to be covered by the GNU General Public
# License. However the source code for this file must still be made available
# in accordance with section (3) of the GNU General Public License.
#
# This exception does not invalidate any other reasons why a work based on
# this file might be covered by the GNU General Public License.
#
# Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
# at http://sources.redhat.com/ecos/ecos-license
# -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Contributors:   gthomas, jskov
# Date:           2001-04-02
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_AMD_PCNET {
    display       "AMD PCNET compatible ethernet driver"
    description   "Ethernet driver for AMD PCNET compatible controllers."

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_IO_ETH_DRIVERS

    active_if     CYGINT_DEVS_ETH_AMD_PCNET_REQUIRED

    include_dir   .
    include_files ; # none _exported_ whatsoever
    compile       -library=libextras.a if_pcnet.c

    define_proc {
        puts $::cdl_header "#include <pkgconf/system.h>";
        puts $::cdl_header "#include CYGDAT_DEVS_ETH_AMD_PCNET_CFG";
    }

    cdl_option CYGNUM_DEVS_ETH_AMD_PCNET_DEV_COUNT {
	display "Number of supported interfaces."
	calculated    { CYGINT_DEVS_ETH_AMD_PCNET_REQUIRED }
        flavor        data
	description   "
	    This option selects the number of PCI ethernet interfaces to
            be supported by the driver."
    }

    cdl_option CYGSEM_DEVS_ETH_AMD_PCNET_FORCE_10MBPS {
        display       "Force negotiation of a 10Mbps link"
        flavor        bool
        default_value 0
        description   "
          If this option is enabled then the driver will force the chipset
          to negotiate only for a 10Mbps link (rather than a 100Mbps
          link)."
    }

    cdl_component CYGPKG_DEVS_ETH_AMD_PCNET_OPTIONS {
        display "PCNET ethernet driver build options"
        flavor  none
	no_define

        cdl_option CYGPKG_DEVS_ETH_AMD_PCNET_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building the PCNET ethernet driver package.
                These flags are used in addition
                to the set of global flags."
        }
    }
}
