# ====================================================================
#
#      ser_mips_ref4955.cdl
#
#      eCos serial MIPS/REF4955 configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  gthomas
# Contributors:
# Date:           2000-05-24
#
#####DESCRIPTIONEND####
#
# ====================================================================


cdl_package CYGPKG_IO_SERIAL_MIPS_REF4955 {
    display       "REF4955 serial device drivers"

    parent        CYGPKG_IO_SERIAL_DEVICES
    active_if     CYGPKG_IO_SERIAL
    active_if     CYGPKG_HAL_MIPS_TX49_REF4955

    requires      CYGPKG_ERROR
    include_dir   cyg/io

    description   "
           This option enables the serial device drivers for the
           REF4955."
    doc           redirect/ecos-device-drivers.html

    # FIXME: This really belongs in the GENERIC_16X5X package
    cdl_interface CYGINT_IO_SERIAL_GENERIC_16X5X_REQUIRED {
        display   "Generic 16x5x serial driver required"
    }

    define_proc {
        puts $::cdl_system_header "/***** serial driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_GENERIC_16X5X_INL <cyg/io/mips_tx49_ref4955_ser.inl>"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_GENERIC_16X5X_CFG <pkgconf/io_serial_mips_ref4955.h>"
        puts $::cdl_system_header "/*****  serial driver proc output end  *****/"
    }

    cdl_component CYGPKG_IO_SERIAL_MIPS_REF4955_SERIAL0 {
        display       "REF4955 serial port 0 driver"
        flavor        bool
        default_value 1
        description   "
            This option includes the serial device driver for the
            REF4955 port 0."

        implements CYGINT_IO_SERIAL_GENERIC_16X5X_REQUIRED
#        implements CYGINT_IO_SERIAL_FLOW_CONTROL_HW
#        implements CYGINT_IO_SERIAL_LINE_STATUS_HW

        cdl_option CYGDAT_IO_SERIAL_MIPS_REF4955_SERIAL0_NAME {
            display       "Device name for the REF4955 serial port 0 driver"
            flavor        data
            default_value {"\"/dev/ser0\""}
            description   "
                This option sets the name of the serial device for the
                REF4955 port 0."
        }

        cdl_option CYGNUM_IO_SERIAL_MIPS_REF4955_SERIAL0_BAUD {
            display       "Baud rate for the REF4955 serial port 0 driver"
            flavor        data
            legal_values  { 1200 2400 4800 9600 14400 19200 38400 57600 115200}
            default_value 38400
            description   "
                This option specifies the default baud rate (speed)
                for the REF4955 port 0."
        }

        cdl_option CYGNUM_IO_SERIAL_MIPS_REF4955_SERIAL0_BUFSIZE {
            display       "Buffer size for the REF4955 serial port 0 driver"
            flavor        data
            legal_values  0 to 8192
            default_value 128
            description   "
                This option specifies the size of the internal buffers
                used for the REF4955 port 0."
        }
    }

    cdl_component CYGPKG_IO_SERIAL_MIPS_REF4955_SERIAL1 {
        display       "REF4955 serial port 1 driver"
        flavor        bool
        default_value 1
        description   "
            This option includes the serial device driver for the
            REF4955 port 1."

        implements CYGINT_IO_SERIAL_GENERIC_16X5X_REQUIRED
#        implements CYGINT_IO_SERIAL_FLOW_CONTROL_HW
#        implements CYGINT_IO_SERIAL_LINE_STATUS_HW

        cdl_option CYGDAT_IO_SERIAL_MIPS_REF4955_SERIAL1_NAME {
            display       "Device name for the REF4955 serial port 1 driver"
            flavor        data
            default_value {"\"/dev/ser1\""}
            description   "
                This option specifies the name of serial device for
                the REF4955 port 1."
        }

        cdl_option CYGNUM_IO_SERIAL_MIPS_REF4955_SERIAL1_BAUD {
            display       "Baud rate for the REF4955 serial port 1 driver"
            flavor        data
            legal_values  { 1200 2400 4800 9600 14400 19200 38400 57600 115200}
            default_value 38400
            description   "
                This option specifies the default baud rate (speed)
                for the REF4955 port 1."
        }

        cdl_option CYGNUM_IO_SERIAL_MIPS_REF4955_SERIAL1_BUFSIZE {
            display       "Buffer size for the REF4955 serial port 1 driver"
            flavor        data
            legal_values  0 to 8192
            default_value 128
            description   "
                This option specifies the size of the internal buffers
                used for the REF4955 port 1."
        }
    }


    cdl_component CYGPKG_IO_SERIAL_MIPS_REF4955_TESTING {
        display    "Testing parameters"
        flavor     bool
        calculated 1
        active_if  CYGPKG_IO_SERIAL_MIPS_REF4955_SERIAL0
        
        cdl_option CYGPRI_SER_TEST_SER_DEV {
            display       "Serial device used for testing"
            flavor        data
            default_value { CYGDAT_IO_SERIAL_MIPS_REF4955_SERIAL0_NAME }
        }

        define_proc {
            puts $::cdl_header "#define CYGPRI_SER_TEST_CRASH_ID \"ref4955\""
            puts $::cdl_header "#define CYGPRI_SER_TEST_TTY_DEV  \"/dev/tty0\""
        }
    }
}

# EOF ser_mips_ref4955.cdl
