# ====================================================================
#
#      usbs.cdl
#
#      USB slave-side support
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 2000, 2001 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      bartv
# Original data:  bartv
# Contributors:
# Date:           2000-10-04
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_IO_USB_SLAVE {
    display     "USB slave-side support"
    parent      CYGPKG_IO_USB
    include_dir "cyg/io/usb"
    active_if   CYGHWR_IO_USB_SLAVE
    doc         io-usb-slave.html
    
    compile usbs.c

    cdl_interface CYGINT_IO_USB_SLAVE_CLIENTS {
	display         "Number of clients of USB devices"
	description "
	    This counter keeps track of the number of clients of
	    USB devices, especially application-class packages such
	    as the USB-ethernet support. It can be used by USB
	    device drivers for default settings.
	"
    }

    cdl_option CYGGLO_IO_USB_SLAVE_APPLICATION {
	display         "Application code uses USB devices"
	default_value   0
	implements      CYGINT_IO_USB_SLAVE_CLIENTS
	description "
	    If the USB devices are accessed by application code
	    rather than by other packages then enabling this
	    option will cause the USB device drivers to be enabled. 
	"
    }
    
    cdl_option CYGGLO_IO_USB_SLAVE_PROVIDE_DEVTAB_ENTRIES {
	display         "Provide devtab entries by default"
	default_value   CYGPKG_IO
	requires        CYGPKG_IO
	description "
	    The USB slave-side endpoints can typically be accessed in two
	    different ways. There is support for the traditional way of
	    doing I/O with open/read/write calls, which involves the
	    use of devtab entries. It is also possible to use a
	    USB-specific API, defined largely in terms of asynchronous
	    operations and callbacks (the read/write implementation uses
	    these lower-level calls). If neither the application nor
	    any other USB-related packages require the higher-level
            read/write calls then it is possible to save some memory
	    by eliminating the devtab entries.
	"
    }
    
    cdl_interface CYGHWR_IO_USB_SLAVE_OUT_ENDPOINTS {
	display "Number of available host->slave endpoints"
    }
    cdl_interface CYGHWR_IO_USB_SLAVE_IN_ENDPOINTS {
	display "Number of available slave->host endpoints"
    }
}
