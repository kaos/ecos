# ====================================================================
#
#      hal_arm_pid.cdl
#
#      PID board HAL package configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      bartv
# Original data:  gthomas
# Contributors:
# Date:           1999-06-13
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_ARM_PID {
    display       "ARM PID evaluation board"
    parent        CYGPKG_HAL_ARM
    define_header hal_arm_pid.h
    include_dir   cyg/hal
    hardware
    description   "
        The pid HAL package provides the support needed to run
        eCos on an ARM PID evaluation board."

    compile       hal_diag.c pid_misc.c

    implements    CYGINT_HAL_DEBUG_GDB_STUBS
    implements    CYGINT_HAL_DEBUG_GDB_STUBS_BREAK
    implements    CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H   <pkgconf/hal_arm.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_arm_pid.h>"
        puts $::cdl_header ""
        puts $::cdl_header "#define HAL_PLATFORM_CPU    \"ARM 7TDMI\""
        puts $::cdl_header "#define HAL_PLATFORM_BOARD  \"PID\""
        puts $::cdl_header "#define HAL_PLATFORM_EXTRA  \"\""
        puts $::cdl_header ""
    }


    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        legal_values  {"RAM" "ROM"}
        default_value {"RAM"}
	no_define
	define -file system.h CYG_HAL_STARTUP
        description   "
            When targetting the PID eval board it is possible to build
            the system for either RAM bootstrap or ROM bootstrap(s). Select
            'ram' when building programs to load into RAM using onboard
            debug software such as Angel or eCos GDB stubs.  Select 'rom'
            when building a stand-alone application which will be put
            into ROM."

    }

    cdl_option CYGHWR_HAL_ARM_PID_DIAG_PORT {
        display       "Diagnostic serial port"
        flavor        data
        legal_values  0 1
        default_value 0
        description   "
            The PID board has two separate serial ports.  This option
            chooses which of these ports will be used."
    }

    cdl_option CYGHWR_HAL_ARM_PID_DIAG_BAUD {
        display       "Diagnostic serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 115200
        default_value 38400
        description   "
            This option selects the baud rate used for the diagnostic port.
            Note: this should match the value chosen for the GDB port if the
            diagnostic and GDB port are the same."
    }

    cdl_option CYGHWR_HAL_ARM_PID_GDB_PORT {
        display       "GDB serial port"
        flavor        data
        legal_values  0 1
        default_value 0
        description   "
            The PID board has two separate serial ports.  This option
            chooses which of these ports will be used to connect to a host
            running GDB."
    }

    cdl_option CYGHWR_HAL_ARM_PID_GDB_BAUD {
        display       "GDB serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 115200
        default_value 38400
        description   "
            This option controls the baud rate used for the GDB connection."
    }

    cdl_option CYGHWR_HAL_ARM_PID_DIAG_LEDS {
        display          "Enable use of PPx LEDs"
        default_value    0
        description      "
            The PID board has four LEDs labelled PP0-PP3. These can be
            controlled by eCos if jumpers 9-16 on LK11 are
            shorted. Note that this prevents the parallel port from
            being used. See the PID board manual for details.
            
            Enabling this option causes eCos to flash the LEDs during
            early board initialization. See vectors.S for
            details. Before calling cyg_start, PP0 is switched on,
            PP1-3 are switched off. The application code can use the
            function hal_diag_led() to control the LEDs after this
            point."
   }


    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
        display      "Number of communication channels on the board"
        flavor       data
        calculated   2
    }
 
    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
        display          "Debug serial port"
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    CYGHWR_HAL_ARM_PID_GDB_PORT
        description      "
            The PID board has only one serial port. This option
            chooses which port will be used to connect to a host
            running GDB."
     }
 
     cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
         display          "Diagnostic serial port"
         flavor data
         legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
         default_value    CYGHWR_HAL_ARM_PID_DIAG_PORT
         description      "
            The PID board has only one serial port.  This option
            chooses which port will be used for diagnostic output."
     }

    # Real-time clock/counter specifics
    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants"
        flavor        none
    
        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            calculated    1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            calculated    100
        }
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
           calculated    12500
        }
    }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        parent  CYGPKG_NONE
        description   "
	    Global build options including control over
	    compiler flags, linker flags and choice of toolchain."


        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { CYGHWR_THUMB ? "thumb-elf" : "arm-elf" }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { (CYGHWR_THUMB && CYGHWR_HAL_ARM_BIGENDIAN) ? "-mthumb-interwork -mbig-endian -Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority" :
            CYGHWR_THUMB ? "-mthumb-interwork -Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority" :
            (CYGHWR_HAL_ARM_CPU_FAMILY == "ARM9") && CYGHWR_HAL_ARM_BIGENDIAN ? "-mcpu=arm9 -mbig-endian -Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority" :
            (CYGHWR_HAL_ARM_CPU_FAMILY == "ARM9") && ! CYGHWR_HAL_ARM_BIGENDIAN ? "-mcpu=arm9 -Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority" :
            (CYGHWR_HAL_ARM_CPU_FAMILY != "ARM9") && CYGHWR_HAL_ARM_BIGENDIAN ? "-mcpu=arm7tdmi -mbig-endian -Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority" :
            "-mcpu=arm7tdmi -Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority" }
            description   "
                This option controls the global compiler flags which are used to
                compile all packages by default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { (CYGHWR_THUMB && CYGHWR_HAL_ARM_BIGENDIAN) ? "-mthumb-interwork -mbig-endian -g -nostdlib -Wl,--gc-sections -Wl,-static" :
            CYGHWR_THUMB ? "-mthumb-interwork -g -nostdlib -Wl,--gc-sections -Wl,-static" :
            (CYGHWR_HAL_ARM_CPU_FAMILY == "ARM9") && CYGHWR_HAL_ARM_BIGENDIAN ? "-mcpu=arm9 -mbig-endian -g -nostdlib -Wl,--gc-sections -Wl,-static" :
            (CYGHWR_HAL_ARM_CPU_FAMILY == "ARM9") && ! CYGHWR_HAL_ARM_BIGENDIAN ? "-mcpu=arm9 -g -nostdlib -Wl,--gc-sections -Wl,-static" :
            (CYGHWR_HAL_ARM_CPU_FAMILY != "ARM9") && CYGHWR_HAL_ARM_BIGENDIAN ? "-mcpu=arm7tdmi -mbig-endian -g -nostdlib -Wl,--gc-sections -Wl,-static" :
            "-mcpu=arm7tdmi -g -nostdlib -Wl,--gc-sections -Wl,-static" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }

        cdl_option CYGBLD_BUILD_GDB_STUBS {
            display "Build GDB stub ROM image"
            default_value 0
            requires CYGBLD_BUILD_COMMON_GDB_STUBS
            requires { CYG_HAL_STARTUP == "ROM" }
            requires CYGSEM_HAL_ROM_MONITOR
            requires CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT
            requires CYGDBG_HAL_DEBUG_GDB_THREAD_SUPPORT
            requires ! CYGDBG_HAL_COMMON_INTERRUPTS_SAVE_MINIMUM_CONTEXT
            requires ! CYGDBG_HAL_COMMON_CONTEXT_SAVE_MINIMUM
            no_define
            description "
                This option enables the building of the GDB stubs for the
                board. The address of the ELF headers in the image are
                adjusted to ensure loading at an address in memory used
                by the flash tool."

            make -priority 320 {
                <PREFIX>/bin/gdb_module.bin : <PREFIX>/bin/gdb_module.img
                @mv $< $(<:.img=.elf)
                $(OBJCOPY) --strip-debug --change-addresses=0xFC060000 $(<:.img=.elf) $<
                $(OBJCOPY) -O binary $(<:.img=.elf) $@
            }
        }

        cdl_option CYGBLD_BUILD_FLASH_TOOL {
            display "Build flash programming tool"
            default_value 0
            requires { CYG_HAL_STARTUP == "RAM" }
            requires CYGHWR_HAL_ARM_PID_DIAG_PORT == 1
            requires CYGPKG_LIBC
            requires CYGPKG_KERNEL
            no_define
            description "This option enables the building of the flash programming tool for copying the GDB stubs into flash memory."
            make -priority 320 {
                <PREFIX>/bin/prog_flash.img : <PACKAGE>/src/prog_flash.c
                @sh -c "mkdir -p src $(dir $@)"
                $(CC) -c $(INCLUDE_PATH) -Wp,-MD,deps.tmp -I$(dir $<) $(CFLAGS) -o src/prog_flash.o $<
                @echo $@ ": \\" > $(notdir $@).deps
                @echo $(wildcard $(PREFIX)/lib/*) " \\" >> $(notdir $@).deps
                @tail +2 deps.tmp >> $(notdir $@).deps
                @echo >> $(notdir $@).deps
                @rm deps.tmp
                $(CC) $(LDFLAGS) -L$(PREFIX)/lib -Ttarget.ld -o $@ src/prog_flash.o
            }
        }

        cdl_option CYGBLD_BUILD_FLASH_TOOL_BE {
            display "Build flash programming tool for BE images on LE boards"
            default_value 0
            requires { CYG_HAL_STARTUP == "RAM" }
            requires CYGHWR_HAL_ARM_PID_DIAG_PORT == 1
            requires CYGPKG_LIBC
            requires CYGPKG_KERNEL
            no_define
            description "This option enables the building of the flash
                         programming tool for copying the GDB stubs
                         into flash memory. The tool built by enabling
                         this option must be used when programming BE
                         images on LE boards."
            make -priority 320 {
                <PREFIX>/bin/prog_flash_BE_image_LE_system.img : <PACKAGE>/src/prog_flash.c
                @sh -c "mkdir -p src $(dir $@)"
                $(CC) -DBE_IMAGE -c $(INCLUDE_PATH) -Wp,-MD,deps.tmp -I$(dir $<) $(CFLAGS) -o src/prog_flash_be.o $<
                @echo $@ ": \\" > $(notdir $@).deps
                @echo $(wildcard $(PREFIX)/lib/*) " \\" >> $(notdir $@).deps
                @tail +2 deps.tmp >> $(notdir $@).deps
                @echo >> $(notdir $@).deps
                @rm deps.tmp
                $(CC) $(LDFLAGS) -L$(PREFIX)/lib -Ttarget.ld -o $@ src/prog_flash_be.o
            }
        }
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { CYG_HAL_STARTUP == "RAM" ? "arm_pid_ram" : \
                                                "arm_pid_rom" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_pid_ram.ldi>" : \
                                                    "<pkgconf/mlt_arm_pid_rom.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_pid_ram.h>" : \
                                                    "<pkgconf/mlt_arm_pid_rom.h>" }
        }
    }


    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "ROM" }
        description   "
            Enable this option if this program is to be used as a ROM monitor,
            i.e. applications will be loaded into RAM on the board, and this
            ROM monitor may process exceptions or interrupts generated from the
            application. This enables features such as utilizing a separate
            interrupt stack when exceptions are generated."
    }

    cdl_component CYGPKG_CYGMON_HAL_OPTIONS {
        display       "CygMon HAL options"
        flavor        none
        no_define
        parent        CYGPKG_CYGMON
        active_if     CYGPKG_CYGMON
        requires      CYGPKG_IO_SERIAL_ARM_PID
        requires      {(CYGDAT_CYGMON_CONSOLE_DEV != "\"/dev/ser0\"") || \
                       (CYGPKG_IO_SERIAL_ARM_PID_SERIAL0 &&              \
                       (CYGNUM_IO_SERIAL_ARM_PID_SERIAL0_BUFSIZE == 512))}
        requires      {(CYGDAT_CYGMON_CONSOLE_DEV != "\"/dev/ser1\"") || \
                       (CYGPKG_IO_SERIAL_ARM_PID_SERIAL1 &&              \
                       (CYGNUM_IO_SERIAL_ARM_PID_SERIAL1_BUFSIZE == 512))}
        description   "
            This option also lists the target's requirements for a valid CygMon
            configuration."


        cdl_option CYGDAT_CYGMON_CONSOLE_DEV {
            display       "Serial port for default console"
            flavor data
            default_value { "\"/dev/ser0\"" }
            description   "
                This option selects the physical device to use as the default
                console device for CygMon."

        }

        cdl_option CYGBLD_BUILD_CYGMON_BIN {
            display       "Build CygMon ROM binary image"
            active_if     CYGBLD_BUILD_CYGMON
            default_value 1
            no_define
            description "This option enables the conversion of the CygMon ELF
                         image to a binary image suitable for ROM programming."
    
            make -priority 325 {
                <PREFIX>/bin/cygmon.bin : <PREFIX>/bin/cygmon.elf
                $(OBJCOPY) --strip-debug --change-addresses=0xFC060000 $< $(@:.bin=.img) 
                $(OBJCOPY) -O srec $< $(@:.bin=.srec)
                $(OBJCOPY) -O binary $< $@
            }
        }
    }

    cdl_option CYGSEM_HAL_USE_ROM_MONITOR {
         display       "Work with a ROM monitor"
         flavor        booldata
         legal_values  { "Generic" "GDB_stubs" }
         default_value { CYG_HAL_STARTUP == "RAM" ? "GDB_stubs" : 0 }
         parent        CYGPKG_HAL_ROM_MONITOR
         requires      { CYG_HAL_STARTUP == "RAM" }
         description   "
             Support can be enabled for different varieties of ROM monitor.
             This support changes various eCos semantics such as the encoding
             of diagnostic output, or the overriding of hardware interrupt
             vectors.
             Firstly there is \"Generic\" support which prevents the HAL
             from overriding the hardware vectors that it does not use, to
             instead allow an installed ROM monitor to handle them. This is
             the most basic support which is likely to be common to most
             implementations of ROM monitor.
             \"GDB_stubs\" provides support when GDB stubs are included in
             the ROM monitor or boot ROM."
     }

}
