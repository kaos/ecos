# ====================================================================
#
#      hal_arm_ebsa285.cdl
#
#      AEB1 board HAL package configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  hmt
# Contributors:
# Date:           1999-08-12
#
#####DESCRIPTIONEND####
#
# ====================================================================
cdl_package CYGPKG_HAL_ARM_EBSA285 {
    display       "Intel EBSA285 StrongARM evaluation boards"
    parent        CYGPKG_HAL_ARM
    define_header hal_arm_ebsa285.h
    include_dir   cyg/hal
    hardware
    description   "
        The EBSA285 HAL package provides the support needed to run
        eCos on a Intel EBSA285 StrongARM eval board."

    compile hal_diag.c plf_stub.c ebsa285_misc.c mem285.S

    implements    CYGINT_HAL_DEBUG_GDB_STUBS
    implements    CYGINT_HAL_DEBUG_GDB_STUBS_BREAK

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H   <pkgconf/hal_arm.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_arm_ebsa285.h>"
    }

    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        default_value {"RAM"}
        legal_values  {"RAM" "ROM"}
	no_define
	define -file system.h CYG_HAL_STARTUP
        description   "
           When targetting the EBSA285 eval board it is possible to build
           the system for either RAM bootstrap or ROM bootstrap(s). Select
           'ram' when building programs to load into RAM using onboard
           debug software such as Angel or eCos GDB stubs.  Select 'rom'
           when building a stand-alone application which will be put
           into ROM.  Selection of 'stubs' is for the special case of
           building the eCos GDB stubs themselves."
   }

   cdl_option CYGHWR_HAL_ARM_EBSA285_PCI_MEM_MAP_BASE {
       display            "Base of memory accessible via PCI space"
       flavor             data
       legal_values       0 to 0x01000000
       default_value      0x00f00000
       active_if          CYGPKG_IO_PCI
       description "
           This option determines the base of the EBSA memory which
           can be accessed via the PCI bus. The default is to allow
           access to the upper 1MB of a 16MB system. Change in 256kB
           increments."
   }

   cdl_option CYGHWR_HAL_ARM_EBSA285_PCI_MEM_MAP_SIZE {
       display            "Size of memory accessible via PCI space"
       flavor             data
       legal_values       0 to 0x01000000
       default_value      0x00100000
       active_if          CYGPKG_IO_PCI
       description "
           This option determines the size of the EBSA memory which
           can be accessed via the PCI bus. The default is to allow
           access to the upper 1MB of a 16MB system. Change in 256kB
           increments."
   }

    # Real-time clock/counter specifics
    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants"
        flavor        none
    
        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            calculated    1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            calculated    100
        }
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
            calculated    36800        ;# Timer3 clock is 3.68MHz
        }
    }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        description   "
	    Global build options including control over
	    compiler flags, linker flags and choice of toolchain."


        parent  CYGPKG_NONE

        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "arm-elf" }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { "-mcpu=strongarm -Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority" }
            description   "
                This option controls the global compiler flags which are used to
                compile all packages by default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { "-Wl,--gc-sections -Wl,-static -g -O2 -nostdlib" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }

        cdl_option CYGBLD_BUILD_GDB_STUBS {
            display "Build GDB stub ROM image"
            default_value 0
            requires { CYG_HAL_STARTUP == "ROM" }
            requires CYGSEM_HAL_ROM_MONITOR
            requires CYGBLD_BUILD_COMMON_GDB_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
            requires ! CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT
            requires ! CYGDBG_HAL_DEBUG_GDB_THREAD_SUPPORT
            requires ! CYGDBG_HAL_COMMON_INTERRUPTS_SAVE_MINIMUM_CONTEXT
            requires ! CYGDBG_HAL_COMMON_CONTEXT_SAVE_MINIMUM
            no_define
            description "
                This option enables the building of the GDB stubs for the
                board. The common HAL controls takes care of most of the
                build process, but the final conversion from ELF image to
                binary data is handled by the platform CDL, allowing
                relocation of the data if necessary."

            make -priority 320 {
                <PREFIX>/bin/gdb_module.bin : <PREFIX>/bin/gdb_module.img
                $(OBJCOPY) -O binary $< $@
            }
        }
    }

    cdl_component CYGPKG_HAL_ARM_EBSA285_OPTIONS {
        display "StrongARM EBSA285 build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_HAL_ARM_EBSA285_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the StrongARM EBSA285 HAL. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_HAL_ARM_EBSA285_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the StrongARM EBSA285 HAL. These flags are removed from
                the set of global flags if present."
        }

        cdl_option CYGPKG_HAL_ARM_EBSA285_TESTS {
            display "StrongARM EBSA285 tests"
            flavor  data
            no_define
            calculated { "tests/sdram0" }
            description   "
                This option specifies the set of tests for the StrongARM EBSA285 HAL."
        }
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { CYG_HAL_STARTUP == "RAM" ? "arm_ebsa285_ram" : \
	                                        "arm_ebsa285_rom" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_ebsa285_ram.ldi>" : \
                                                    "<pkgconf/mlt_arm_ebsa285_rom.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_ebsa285_ram.h>" : \
                                                    "<pkgconf/mlt_arm_ebsa285_rom.h>" }
        }
    }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "ROM" }
        description   "
            Enable this option if this program is to be used as a ROM monitor,
            i.e. applications will be loaded into RAM on the board, and this
            ROM monitor may process exceptions or interrupts generated from the
            application. This enables features such as utilizing a separate
            interrupt stack when exceptions are generated."
    }
}
