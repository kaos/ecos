# ====================================================================
#
#	intel_i82559_eth_drivers.cdl
#
#	Intel 82559 ethernet driver
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      hmt
# Original data:  hmt
# Contributors:	  hmt, gthomas, jskov
# Date:           2000-02-01
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_INTEL_I82559 {
    display       "Intel 82559 ethernet driver"
    description   "Ethernet driver for Intel 82559 controller."

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if     CYGPKG_IO_ETH_DRIVERS

    active_if     CYGINT_DEVS_ETH_INTEL_I82559_REQUIRED
    implements    CYGINT_IO_ETH_MULTICAST

    include_dir   cyg/devs/eth

    # SNMP demands to know stuff; this sadly makes us break the neat
    # abstraction of the device having nothing exported.
    include_files include/i82559_info.h
    # and tell them that it is available
    define_proc {
	puts $::cdl_system_header \
       "#define CYGBLD_DEVS_ETH_DEVICE_H <pkgconf/devs_eth_intel_i82559.h>"

        puts $::cdl_header "#include CYGDAT_DEVS_ETH_INTEL_I82559_CFG";
    }

    compile       -library=libextras.a if_i82559.c

    cdl_option CYGDBG_DEVS_ETH_INTEL_I82559_CHATTER {
	display "Prints ethernet device status info during startup"
	default_value 0
	description   "
	    The ethernet device initialization code can print lots of info
	    to confirm that it has found the devices on the PCI bus, read
	    the MAC address from EEPROM correctly, and so on, and also
	    displays the mode (10/100MHz, half/full duplex) of the
	    connection."
    }

    cdl_option CYGNUM_DEVS_ETH_INTEL_I82559_DEV_COUNT {
	display "Number of supported interfaces."
	calculated    { CYGINT_DEVS_ETH_INTEL_I82559_REQUIRED }
        flavor        data
	description   "
	    This option selects the number of PCI ethernet interfaces to
            be supported by the driver."
    }

    cdl_component CYGDBG_DEVS_ETH_INTEL_I82559_KEEP_STATISTICS {
	display "Keep Ethernet statistics"
	default_value 1
	description   "
	    The ethernet device can maintain statistics about the network,
	    specifically a great variety of error rates which are useful
	    for network management.  SNMP for example uses this
	    information.  There is some performance cost in maintaining
	    this information; disable this option to recoup that."

	cdl_option CYGDBG_DEVS_ETH_INTEL_I82559_KEEP_82559_STATISTICS {
	    display "Keep i82559 Internal statistics"
	    default_value 1
	    description   "
	        The i82559 keeps internal counters, and it is possible to
	        acquire these.  But the i82559 (reputedly) does not service
	        the network whilst uploading the data to RAM from its
	        internal registers.  If throughput is a problem, disable
	        this option to acquire only those statistics gathered by
	        software, so that the i82559 never sleeps."
	}
    }

    cdl_component CYGPKG_DEVS_ETH_INTEL_I82559_WRITE_EEPROM {
	display "SIOCSIFHWADDR records MAC address in EEPROM"
	default_value 0
	description   "
	    The ioctl() socket call with operand SIOCSIFHWADDR sets the
	    interface hardware address - the MAC address or ethernet
	    address.  This option causes the new MAC address to be written
	    into the EEPROM associated with the interface, so that the new
	    MAC address is permanently recorded.  Doing this should be a
	    carefully chosen decision, hence this option."
    }

    cdl_option CYGNUM_DEVS_ETH_INTEL_I82559_MAX_RX_DESCRIPTORS {
        display       "Maximum number of RX descriptors"
        flavor  data
        default_value { CYGPKG_REDBOOT ? 4 : 128 }
        define        MAX_RX_DESCRIPTORS
        description   "
                An RX descriptor is used for each ethernet frame required
                to be passed to the upper networking layers. This option
                sets the maximum number of these. Higher numbers use more
                memory, lower numbers will reduce performance. The system
                appears to work OK with as few as 8 descriptors but limps
                painfully with only 4. Performance is better with more than
                8, but assuming the size of non-cached (so useless for anything
                else) memory window is 1Mb, we might as well use it all.
                128 RX and TX descriptors uses the whole 1Mb, near enough."
    }
    
    cdl_option CYGNUM_DEVS_ETH_INTEL_I82559_MAX_TX_DESCRIPTORS {
        display       "Maximum number of TX descriptors"
        flavor  data
        default_value { CYGPKG_REDBOOT ? 4 : 128 }
        define        MAX_TX_DESCRIPTORS
        description   "
                A TX descriptor is used for each ethernet frame passed down
                from upper networking layers for transmission. This option
                sets the maximum number of these. Higher numbers use more
                memory, lower numbers will reduce performance. The system
                appears to work OK with as few as 8 descriptors but limps
                painfully with only 4. Performance is better with more than
                8, but assuming the size of non-cached (so useless for anything
                else) memory window is 1Mb, we might as well use it all.
                128 RX and TX descriptors uses the whole 1Mb, near enough."
    }

    cdl_component CYGPKG_DEVS_ETH_INTEL_I82559_OPTIONS {
        display "Intel 82559 ethernet driver build options"
        flavor  none
	no_define

        cdl_option CYGPKG_DEVS_ETH_INTEL_I82559_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building the Intel 82559 ethernet driver
                package. These flags are used in addition to the set of
                global flags."
        }
    }
}
# EOF intel_i82559_eth_drivers.cdl
