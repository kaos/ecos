# ====================================================================
#
#      hal_v85x_v850.cdl
#
#      NEC/V850 variant architectural HAL package configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Contributors:
# Date:           2000-03-09
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_V85X_V850 {
    display       "V850 variant"
    parent        CYGPKG_HAL_V85X
    implements    CYGINT_HAL_V85X_VARIANT
    hardware
    include_dir   cyg/hal
    define_header hal_v85x_v850.h
    description   "
           The V850 variant HAL package provides generic support
           for this processor architecture. It is also necessary to
           select a specific target platform HAL package."

    define_proc {
        puts $::cdl_header "#include <pkgconf/hal_v85x.h>"
    }

    compile v850_stub.c v850_misc.c context.S

    cdl_interface CYGINT_HAL_V85X_VARIANT_SA1 {
        display  "Defined if CPU is a V850/SA1"
    }

    cdl_interface CYGINT_HAL_V85X_VARIANT_SB1 {
        display  "Defined if CPU is a V850/SB1"
    }

    make {
        <PREFIX>/lib/target.ld: <PACKAGE>/src/v85x_v850.ld
        $(CC) -E -P -Wp,-MD,target.tmp -DEXTRAS=1 -xc $(INCLUDE_PATH) $(CFLAGS) -o $@ $<
        @echo $@ ": \\" > $(notdir $@).deps
        @tail +2 target.tmp >> $(notdir $@).deps
        @echo >> $(notdir $@).deps
        @rm target.tmp
    }

    cdl_option CYGBLD_LINKER_SCRIPT {
        display "Linker script"
        flavor data
	no_define
        calculated  { "src/v85x_v850.ld" }
    }

}
