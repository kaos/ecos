# ====================================================================
#
#      ser_sparclite_sleb.cdl
#
#      eCos serial SPARClite/SLEB configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  gthomas
# Contributors:
# Date:           1999-07-14
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_IO_SERIAL_SPARCLITE_SLEB {
    display       "SPARClite SLEB serial device drivers"

    parent        CYGPKG_IO_SERIAL_DEVICES
    active_if     CYGPKG_IO_SERIAL
    active_if     CYGPKG_HAL_SPARCLITE_SLEB

    requires      CYGPKG_ERROR
    include_dir   cyg/io
    include_files ; # none _exported_ whatsoever
    description   "
           This option enables the serial device drivers for the
           SPARClite SLEB."
    doc           redirect/ecos-device-drivers.html

    compile       -library=libextras.a   sleb_sdtr.c

    define_proc {
        puts $::cdl_system_header "/***** serial driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_DEVICE_HEADER <pkgconf/io_serial_sparclite_sleb.h>"
        puts $::cdl_system_header "/*****  serial driver proc output end  *****/"
    }

cdl_component CYGPKG_IO_SERIAL_SPARCLITE_SLEB_CON1 {
    display       "SPARClite SLEB serial CON1 port driver"
    flavor        bool
    default_value 1
    description   "
        This option includes the serial device driver for the SPARClite
        SLEB CON1 port."

    cdl_option CYGDAT_IO_SERIAL_SPARCLITE_SLEB_CON1_NAME {
        display       "Device name for SPARClite SLEB serial CON1 port"
        flavor        data
        default_value {"\"/dev/ser0\""}
        description   "
            This option specifies the device name for the SPARClite SLEB
            CON1 port."
    }

    cdl_option CYGNUM_IO_SERIAL_SPARCLITE_SLEB_CON1_BAUD {
        display       "Baud rate for the SPARClite SLEB serial CON1 driver"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                        4800 7200 9600 14400 19200 38400 57600 115200 230400
        }
        default_value 19200
        description   "
            This option specifies the default baud rate (speed) for the
            SPARClite SLEB CON1."
    }

    cdl_option CYGNUM_IO_SERIAL_SPARCLITE_SLEB_CON1_BUFSIZE {
        display       "Buffer size for the SPARClite SLEB serial CON1 driver"
        flavor        data
        legal_values  0 to 8192
        default_value 128
        description   "
            This option specifies the size of the internal buffers used for
            the SPARClite SLEB CON1."
    }
}
cdl_component CYGPKG_IO_SERIAL_SPARCLITE_SLEB_CON2 {
    display       "SPARClite SLEB serial CON2 port driver"
    flavor        bool
    default_value 1
    description   "
        This option includes the serial device driver for the SPARClite 
        SLEB CON2 port."

    cdl_option CYGDAT_IO_SERIAL_SPARCLITE_SLEB_CON2_NAME {
        display       "Device name for SPARClite SLEB serial CON2 port"
        flavor        data
        default_value {"\"/dev/ser1\""}
        description   "
            This option specifies the device name for the SPARClite SLEB
            CON2 port."
    }

    cdl_option CYGNUM_IO_SERIAL_SPARCLITE_SLEB_CON2_BAUD {
        display       "Baud rate for the SPARClite SLEB serial CON2 driver"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 230400
        }
        default_value 19200
        description   "
            This option specifies the default baud rate (speed) for the
            SPARClite SLEB CON2."
    }

    cdl_option CYGNUM_IO_SERIAL_SPARCLITE_SLEB_CON2_BUFSIZE {
        display       "Buffer size for the SPARClite SLEB serial CON2 driver"
        flavor        data
        legal_values  0 to 8192
        default_value 128
        description   "
            This option specifies the size of the internal buffers used for 
            the SPARClite SLEB CON2."
    }
}

    cdl_component CYGPKG_IO_SERIAL_SPARCLITE_SLEB_OPTIONS {
        display "Serial device driver build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_IO_SERIAL_SPARCLITE_SLEB_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_IO_SERIAL_SPARCLITE_SLEB_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are removed from
                the set of global flags if present."
        }
    }

    cdl_component CYGPKG_IO_SERIAL_SPARCLITE_SLEB_TESTING {
        display    "Testing parameters"
        flavor     bool
        calculated 1
        active_if  CYGPKG_IO_SERIAL_SPARCLITE_SLEB_CON1

        implements CYGINT_IO_SERIAL_TEST_SKIP_38400
        implements CYGINT_IO_SERIAL_TEST_SKIP_57600
        implements CYGINT_IO_SERIAL_TEST_SKIP_115200

        cdl_option CYGPRI_SER_TEST_SER_DEV {
            display       "Serial device used for testing"
            flavor        data
            default_value { CYGDAT_IO_SERIAL_SPARCLITE_SLEB_CON1_NAME }
        }

        define_proc {
            puts $::cdl_header "#define CYGPRI_SER_TEST_CRASH_ID \"sparcl\""
            puts $::cdl_header "#define CYGPRI_SER_TEST_TTY_DEV  \"/dev/tty0\""
            puts $::cdl_header "#define CYGPRI_SER_TEST_OVERRIDE_INT_1 CYGNUM_HAL_INTERRUPT_9"
            puts $::cdl_header "#define CYGPRI_SER_TEST_OVERRIDE_INT_2 CYGNUM_HAL_INTERRUPT_10"
        }
    }
}

# EOF ser_sparclite_sleb.cdl
