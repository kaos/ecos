# ====================================================================
#
#      hal_powerpc.cdl
#
#      PowerPC architectural HAL package configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  bartv
# Contributors:
# Date:           1999-11-02
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_POWERPC {
    display  "PowerPC architecture"
    parent        CYGPKG_HAL
    hardware
    include_dir   cyg/hal
    define_header hal_powerpc.h
    description   "
        The PowerPC architecture HAL package provides generic
        support for this processor architecture. It is also
        necessary to select a specific target platform HAL
        package."

    cdl_interface CYGINT_HAL_POWERPC_VARIANT {
        display  "Number of variant implementations in this configuration"
        requires 1 == CYGINT_HAL_POWERPC_VARIANT
    }

    compile       hal_misc.c context.S ppc_stub.c hal_intr.c

    # The "-o file" is a workaround for CR100958 - without it the
    # output file would end up in the source directory under CygWin.
    # n.b. grep does not behave itself under win32
    make -priority 1 {
        <PREFIX>/include/cyg/hal/ppc_offsets.inc : <PACKAGE>/src/hal_mk_defs.c
        $(CC) $(CFLAGS) $(INCLUDE_PATH) -Wp,-MD,ppc_offsets.tmp -o hal_mk_defs.tmp -S $<
        fgrep .equ hal_mk_defs.tmp | sed s/#// > $@
        @echo $@ ": \\" > $(notdir $@).deps
        @tail +2 ppc_offsets.tmp >> $(notdir $@).deps
        @echo >> $(notdir $@).deps
        @rm ppc_offsets.tmp hal_mk_defs.tmp
    }

    make {
        <PREFIX>/lib/vectors.o : <PACKAGE>/src/vectors.S
        $(CC) -Wp,-MD,vectors.tmp $(INCLUDE_PATH) $(CFLAGS) -c -o $@ $<
        @echo $@ ": \\" > $(notdir $@).deps
        @tail +2 vectors.tmp >> $(notdir $@).deps
        @echo >> $(notdir $@).deps
        @rm vectors.tmp
    }

    make {
        <PREFIX>/lib/target.ld: <PACKAGE>/src/powerpc.ld
        $(CC) -E -P -Wp,-MD,target.tmp -DEXTRAS=1 -xc $(INCLUDE_PATH) $(CFLAGS) -o $@ $<
        @echo $@ ": \\" > $(notdir $@).deps
        @tail +2 target.tmp >> $(notdir $@).deps
        @echo >> $(notdir $@).deps
        @rm target.tmp
    }


    cdl_option CYGSEM_HAL_POWERPC_COPY_VECTORS {
        display       "Copy exception vectors to RAM"
        default_value { (CYG_HAL_STARTUP != "RAM" ||
                         CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS) ? 1 : 0 }
        requires      ! CYGSEM_HAL_USE_ROM_MONITOR
        description   "
            Enable this option to force exception vectors to be copied
            to address 0 on startup. For RAM startup this is normally
            disabled since the vectors would already have been provided
            by the GDB stubs - but it's possible to override, thus taking
            full control of the target. For ROM startup it is desirable to
            enable this option for performance reasons (accessing vectors
            in ROM is normally slower) - but if memory is tight the vectors
            can be left in ROM."
    }

    cdl_option CYGDBG_HAL_POWERPC_FRAME_WALLS {
        display       "Exception stack-frame walls"
        default_value 0
        description   "
            Enable this option to put \"walls\" around the exception
            frames. This can ease analyzing the stack contents when
            debugging."
    }

    cdl_component CYGPKG_HAL_POWERPC_OPTIONS {
        display "PowerPC build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_HAL_POWERPC_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the PowerPC HAL. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_HAL_POWERPC_CFLAGS_REMOVE {
            display "Supressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the PowerPC HAL. These flags are removed from
                the set of global flags if present."
        }

        cdl_option CYGPKG_HAL_POWERPC_TESTS {
            display "PowerPC tests"
            flavor  data
            no_define
            calculated { "" }
            description   "
                This option specifies the set of tests for the PowerPC HAL."
        }
    }

    cdl_option CYGBLD_LINKER_SCRIPT {
        display "Linker script"
        flavor data
	no_define
        calculated  { "src/powerpc.ld" }
    }
}
