# ====================================================================
#
#      hal_arm_lpc24xx.cdl
#
#      NXP LPC24XX HAL package configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
## Copyright (C) 2003 Nick Garnett <nickg@calivar.com>
## Copyright (C) 2004 eCosCentric Limited 
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Uwe Kindler
# Contributors:   gthomas, tkoeller, tdrury, nickg
# Date:           2008-07-05
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_ARM_LPC24XX {
    display       "NXP LPC24XX variant HAL"
    parent        CYGPKG_HAL_ARM
    define_header hal_arm_lpc24xx.h
    include_dir   cyg/hal
    hardware
    description   "
        The LPC24XX HAL package provides the support needed to run
        eCos on NXP LPC24XX based targets."

    compile       hal_diag.c lpc24xx_misc.c

    implements    CYGINT_HAL_DEBUG_GDB_STUBS
    implements    CYGINT_HAL_DEBUG_GDB_STUBS_BREAK
    implements    CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT
    implements    CYGINT_HAL_VIRTUAL_VECTOR_COMM_BAUD_SUPPORT
    implements    CYGINT_HAL_ARM_ARCH_ARM7
    implements    CYGINT_HAL_ARM_THUMB_ARCH

    # Let the architectural HAL see this variant's files
    define_proc {
        puts $::cdl_header "#define CYGBLD_HAL_VAR_INTS_H <cyg/hal/hal_var_ints.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_ARM_VAR_IO_H"
        puts $::cdl_system_header "#define CYGBLD_HAL_ARM_VAR_ARCH_H"
    }

    cdl_component CYGHWR_HAL_ARM_LPC24XX {
        display        "LPC24XX variant used"
        flavor         data
        default_value  { "LPC246x" }
        legal_values   { "LPC246x" "LPC2458" "LPC2460" "LPC2468" "LPC2470" 
                         "LPC2478"}
        description    "
             The LPC24XX microcontroller family has several variants,
             the main differences being the amount of on-chip RAM,
             flash and peripherals. This option allows the platform
             HALs to select the specific microcontroller being used."

        cdl_option CYGHWR_HAL_ARM_LPC24XX_FAMILY {
            display       "LPC24XX variant family"
            flavor        data
            calculated    {
                is_substr(CYGHWR_HAL_ARM_LPC24XX, "LPC246") ? 
                   "LPC246X" : "LPC24XX"
                          }
            description   "
                This specifies the family that the processor
                belongs to. This is useful as it defines certain common
                characteristics which affect which features should be
                available in the HAL."
        }
    }
    
    # This is going to get really messy before long as the number of parts
    # explodes. Its useful to know the actual part in use, but its just as
    # useful to know which family it belongs to. LPC210x shouldn't really
    # be in the list of devices, but will probably break something if removed.
    cdl_component CYGHWR_HAL_ARM_LPC2XXX {
        display        "LPC2XXX variant used"
        flavor         data
        calculated     CYGHWR_HAL_ARM_LPC24XX
        description    "
             This option is only here for compatibility reasons because some of
             the LPC2XXX device drivers rely on these definitions. If this
             is defined here, the LPC24XX variant can use the LPC2XXX device
             drivers for on-chip peripherals."

        cdl_option CYGHWR_HAL_ARM_LPC2XXX_FAMILY {
            display       "LPC2XXX variant family"
            flavor        data
            calculated    CYGHWR_HAL_ARM_LPC24XX_FAMILY
            description   "
                 This option is only here for compatibility reasons
                 because some of the LPC2XXX device drivers rely on
                 these definitions. If this is defined here, the
                 LPC24XX variant can use the LPC2XXX device drivers
                 for on-chip peripherals."
        }
        
        cdl_option CYGHWR_HAL_ARM_LPC2XXX_VARIANT_VERSION {
            display       "LPC2XXX variant version"
            flavor        data
            calculated    {
                is_substr(CYGHWR_HAL_ARM_LPC2XXX, "LPC21") ? 1 :
                is_substr(CYGHWR_HAL_ARM_LPC2XXX, "LPC22") ? 2 :
                is_substr(CYGHWR_HAL_ARM_LPC2XXX, "LPC24") ? 4 : 0
                          }
            description   "
                This specifies the variant version that the processor
                belongs to. Some common characteristics may be 
                different in newer LPC2xxx versions. I.e. the LPC24xx variants
                are significant different from former LPC2xxx variants." 
        }
    }

    # Important! Be very careful changing this value. That will always
    # enter the LPC24XX bootloader after reset and consequently will
    # never run your code. You must know what you are doing. Look at
    # arch. vectors.S for details.
    cdl_option CYGNUM_HAL_ARM_VECTOR_0x14 {
        display       "ARM vector at 0x14"
        flavor        data
        default_value 0xB4405F62
        legal_values  0 to 0xFFFFFFFF
        description "
           In order to detect if a valid program is present, every
           user program must have a program signature. This signature
           is a word-wide number that is stored in the unused
           location in the ARM7 vector table at 0x00000014. The
           program signature is the two's compliment of the checksum
           of the ARM vector table."
    }

    cdl_component CYGNUM_HAL_ARM_LPC24XX_CLOCKING {
        display       "Clocking"
        flavor        none

        cdl_option CYGNUM_HAL_ARM_LPC24XX_PLL_MUL {
            display       "PLL multiplier"
            flavor        data
            legal_values  6 to 32767
            default_value { 12 }
        }
    
        cdl_option CYGNUM_HAL_ARM_LPC24XX_PLL_DIV {
            display       "PLL divider"
            flavor         data
            legal_values  1 to 32 
            default_value { 1 }
        }

        cdl_option CYGNUM_HAL_ARM_LPC24XX_PLL_OUTPUT {
            display       "PLL output (MHz)"
            flavor         data
            legal_values   275000000 to 290000000
            calculated {  2 * CYGNUM_HAL_ARM_LPC24XX_PLL_MUL * 
                          CYGNUM_HAL_ARM_LPC24XX_XTAL_FREQ / 
                          CYGNUM_HAL_ARM_LPC24XX_PLL_DIV}
            description "
                Normally the PLL output must be in the range of 275 MHz to 
                550 MHz Because of a chip errata the maximum output of the CCO 
                within the PLL block is limited to 290 MHz."
        }
       
        cdl_component CYGNUM_HAL_ARM_LPC24XX_CLOCK_SPEED {
            display       "CPU clock speed"
            flavor        data
            calculated {  2 * CYGNUM_HAL_ARM_LPC24XX_PLL_MUL * 
                          CYGNUM_HAL_ARM_LPC24XX_XTAL_FREQ / 
                          CYGNUM_HAL_ARM_LPC24XX_PLL_DIV / 
                          CYGNUM_HAL_ARM_LPC24XX_CPU_CLK_DIV}
            description "
                The core CPU clock speed is the PLL output divided by the 
                CPU clock divider" 
                
            cdl_option CYGNUM_HAL_ARM_LPC24XX_CPU_CLK_DIV {
                display       "CPU clock divider"
                flavor        data
                legal_values  6 to 256
                default_value { 6 }
                description "
                    The CPU clock divider controls the division of the PLL 
                    output before it is used by the CPU. When the PLL is 
                    bypassed, the division may be by 1. When the PLL is 
                    running, the output must be divided in order to bring the 
                    CPU clock frequency (CCLK) within operating limits. An 8 
                    bit divider allows a range of options, including slowing 
                    CPU operation to a low rate for temporary power savings 
                    without turning off the PLL. Only even values 
                    (2, 4, 6, ..., 256) are supported and can be used. 
                    Warning: Using an odd value (1, 3, 5, ..., 255) when 
                    setting this option may result in incorrect operation of 
                    the device."
             }    
        }
    
        
        cdl_component CYGNUM_HAL_ARM_LPC24XX_USB_CLOCK_SPEED {
            display       "USB clock speed"
            flavor        data
            calculated {  2 * CYGNUM_HAL_ARM_LPC24XX_PLL_MUL * 
                          CYGNUM_HAL_ARM_LPC24XX_XTAL_FREQ / 
                          CYGNUM_HAL_ARM_LPC24XX_PLL_DIV / 
                          CYGNUM_HAL_ARM_LPC24XX_USB_CLK_DIV}
            description "
                The USB clock speed is the PLL output divided by the 
                USB clock divider" 
                
            cdl_option CYGNUM_HAL_ARM_LPC24XX_USB_CLK_DIV {
                display       "USB clock divider"
                flavor        data
                legal_values  1 to 8
                default_value { 6 }
                description "
                    This divider controls the division of the PLL output before 
                    it is used by the USB block. If the PLL is bypassed, the 
                    division may be by 1. In that case, the PLL input frequency 
                    must be 48 MHz, with a 500 ppm tolerance. When the PLL is 
                    running, the output must be divided in order to bring the 
                    USB clock frequency to 48 MHz with a 50% duty cycle. A 
                    4-bit divider allows obtaining the correct USB clock from 
                    any even multiple of 48 MHz (i.e. any mutliple of 96 MHz) 
                    within the PLL operating range."
            }
        }
        
        cdl_component CYGNUM_HAL_ARM_LPC2XXX_CAN_CLK {
            display       "CAN clock speed"
            flavor        data
            calculated   {  CYGNUM_HAL_ARM_LPC24XX_CLOCK_SPEED / 
                            CYGNUM_HAL_ARM_LPC24XX_CAN_CLK_DIV}
            description "
                The CAN clock speed is the CPU clock output divided by the 
                CAN clock divider" 
                
            cdl_option CYGNUM_HAL_ARM_LPC24XX_CAN_CLK_DIV {
                display       "CAN clock divider"
                flavor        data
                legal_values  { 1 2 4 6 }
                default_value { 1 }
                description "
                    This divider selects the peripheral clock for both CAN 
                    channels. The divider divides the CPU clock to get the 
                    clock for the CAN peripherals."
            }
        }      
    }
    
    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants"
        flavor        none

        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            default_value 1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            default_value 100
        }
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
            default_value { ((CYGNUM_HAL_ARM_LPC24XX_CLOCK_SPEED) / 
                              CYGNUM_HAL_RTC_DENOMINATOR) }
        }
    }

    cdl_option CYGHWR_HAL_ARM_LPC24XX_IDLE_PWRSAVE {
        display       "Stop clock in idle loop to save power"
        flavor        bool
        default_value { is_active(CYGPKG_REDBOOT) ? 0 : 1 }
        description   "
           Select this option when it is desired to save power by
           stopping the processor clock in the idle loop. This is
           controlled by the PCON register. Generally this is a good
           thing, but it may be necessary to disable this when
           debugging via JTAG, as stopping the clock can prevent the
           debugger getting control of the system."
    }
    
    cdl_option CYGNUM_HAL_KERNEL_COUNTERS_CLOCK_ISR_DEFAULT_PRIORITY {
	    display		"Default priority for system clock interrupts"
	    flavor		data
	    legal_values  { 0 to 15 }
        default_value 15
	    description "
            There are 16 priority levels, corresponding to the values 0 through 
            15 decimal, of which 15 is the lowest priority. The reset value of 
            these interrupt priority registers defaults all interrupts to the 
            lowest priority, allowing a single write to elevate the priority 
            of an individual interrupt."
    }

}
