# ====================================================================
#
#      hal_powerpc_cogent.cdl
#
#      PowerPC/Cogent board HAL package configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
## Copyright (C) 2003 Gary Thomas
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  bartv
# Contributors:
# Date:           1999-11-02
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_POWERPC_COGENT {
    display       "Cogent PowerPC evaluation board"
    parent        CYGPKG_HAL_POWERPC
    requires      CYGPKG_HAL_POWERPC_MPC8xx
    define_header hal_powerpc_cogent.h
    include_dir   cyg/hal
    description   "
        The cogent HAL package provides the support needed to run
        eCos on a Cogent board equipped with a PowerPC processor."

    compile       hal_diag.c plf_misc.c cogent.S plf_stub.c

    implements    CYGINT_HAL_DEBUG_GDB_STUBS
    implements    CYGINT_HAL_DEBUG_GDB_STUBS_BREAK
    implements    CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT

    requires      { CYGHWR_HAL_POWERPC_MPC8XX == "823" }

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H   <pkgconf/hal_powerpc_mpc8xx.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_powerpc_cogent.h>"
    }

    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        legal_values  {"RAM" "ROM"}
        default_value {"RAM"}
	no_define
	define -file system.h CYG_HAL_STARTUP
        description   "
           When targetting the cogent board it is possible to build
           the system for either RAM bootstrap or ROM bootstrap. RAM
           bootstrap generally requires that the board
           is equipped with ROMs containing a suitable ROM monitor or
           equivalent software that allows GDB to download the eCos
           application on to the board. The ROM bootstrap typically
           requires that the eCos application be blown into EPROMs or
           equivalent technology."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
        display      "Number of communication channels on the board"
        flavor       data
        calculated   3
        description      "
            Channel 0: Serial A, Channel 1: Serial B, Channel 2: LCD"
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
        display          "Debug serial port"
        flavor data
        legal_values     0 to 1
        default_value    1
        description      "
           The Cogent board has two serial ports. This option
           chooses which port will be used to connect to a host
           running GDB."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
        display          "Diagnostic serial port"
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    1
        description      "
           The Cogent board has two serial ports and an LCD.  This option
           chooses which port will be used for diagnostic output."
    }

    cdl_option CYGHWR_HAL_POWERPC_BOARD_SPEED {
        display          "Development board clock speed (MHz)"
        flavor           data
        default_value    33.330
        description      "
           MPC8xx development boards have various system clock speeds
           depending on the processor fitted.  Select the clock speed
           appropriate for your board so that the system can set the serial
           baud rate correctly, amongst other things."
    }

    # Real-time clock/counter specifics
    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants."
        description   "
            Period is busclock/16/100."
        flavor        none
    
        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            calculated    1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            calculated    100
        }
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
            calculated    { (((CYGHWR_HAL_POWERPC_BOARD_SPEED*1000000)/16)/100) }
        }
    }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        parent  CYGPKG_NONE
        description   "
	    Global build options including control over
	    compiler flags, linker flags and choice of toolchain."


        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "powerpc-eabi" }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { "-msoft-float -mcpu=860 -Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority" }
            description   "
                This option controls the global compiler flags which
                are used to compile all packages by
                default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { "-msoft-float -mcpu=860 -g -nostdlib -Wl,--gc-sections -Wl,-static" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }

        cdl_option CYGBLD_BUILD_GDB_STUBS {
            display "Build GDB stub ROM image"
            default_value 0
            requires { CYG_HAL_STARTUP == "ROM" }
            requires CYGSEM_HAL_ROM_MONITOR
            requires CYGBLD_BUILD_COMMON_GDB_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT
            requires CYGDBG_HAL_DEBUG_GDB_THREAD_SUPPORT
            requires ! CYGDBG_HAL_COMMON_INTERRUPTS_SAVE_MINIMUM_CONTEXT
            requires ! CYGDBG_HAL_COMMON_CONTEXT_SAVE_MINIMUM
            no_define
            description "
                This option enables the building of the GDB stubs for the
                board. The common HAL controls takes care of most of the
                build process, but the final conversion from ELF image to
                binary data is handled by the platform CDL, allowing
                relocation of the data if necessary."

            make -priority 320 {
                <PREFIX>/bin/gdb_module.bin : <PREFIX>/bin/gdb_module.img
                $(OBJCOPY) -O binary $< $@
            }
        }
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { CYG_HAL_STARTUP == "RAM" ? "powerpc_cogent_ram" : \
                                                "powerpc_cogent_rom" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_powerpc_cogent_ram.ldi>" : \
                                                    "<pkgconf/mlt_powerpc_cogent_rom.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_powerpc_cogent_ram.h>" : \
                                                    "<pkgconf/mlt_powerpc_cogent_rom.h>" }
        }
    }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "ROM" }
        description   "
            Enable this option if this program is to be used as a ROM monitor,
            i.e. applications will be loaded into RAM on the board, and this
            ROM monitor may process exceptions or interrupts generated from the
            application. This enables features such as utilizing a separate
            interrupt stack when exceptions are generated."
    }
}
