# ====================================================================
#
#      hal_arm_integrator.cdl
#
#      INTEGRATOR board HAL package configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
# -------------------------------------------
# This file is part of eCos, the Embedded Configurable Operating System.
# Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
#
# eCos is free software; you can redistribute it and/or modify it under
# the terms of the GNU General Public License as published by the Free
# Software Foundation; either version 2 or (at your option) any later version.
#
# eCos is distributed in the hope that it will be useful, but WITHOUT ANY
# WARRANTY; without even the implied warranty of MERCHANTABILITY or
# FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
# for more details.
#
# You should have received a copy of the GNU General Public License along
# with eCos; if not, write to the Free Software Foundation, Inc.,
# 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
#
# As a special exception, if other files instantiate templates or use macros
# or inline functions from this file, or you compile this file and link it
# with other works to produce a work based on this file, this file does not
# by itself cause the resulting work to be covered by the GNU General Public
# License. However the source code for this file must still be made available
# in accordance with section (3) of the GNU General Public License.
#
# This exception does not invalidate any other reasons why a work based on
# this file might be covered by the GNU General Public License.
#
# Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
# at http://sources.redhat.com/ecos/ecos-license
# -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      David A Rusling
# Original data:  gthomas
# Contributors:   Philippe Robin
# Date:           November 7, 2000
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_ARM_INTEGRATOR {
    display       "ARM INTEGRATOR evaluation board"
    parent        CYGPKG_HAL_ARM
    define_header hal_arm_integrator.h
    include_dir   cyg/hal
    hardware
    description   "
        The integrator HAL package provides the support needed to run
        eCos on an ARM INTEGRATOR evaluation board."

    compile       hal_diag.c integrator_misc.c 

    implements    CYGINT_HAL_DEBUG_GDB_STUBS
    implements    CYGINT_HAL_DEBUG_GDB_STUBS_BREAK
    implements    CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H   <pkgconf/hal_arm.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_arm_integrator.h>"
        puts $::cdl_header ""
        puts $::cdl_header "#define HAL_PLATFORM_BOARD  \"INTEGRATOR\""
        puts $::cdl_header "#define HAL_PLATFORM_EXTRA  \"\""
        puts $::cdl_header ""
    }

    cdl_component CYGPKG_HAL_ARM_INTEGRATOR_ARM7 {
	display "ARM 7 specialization"
	active_if  !CYGPKG_HAL_ARM_ARM9
	calculated !CYGPKG_HAL_ARM_ARM9

	implements    CYGINT_HAL_ARM_ARCH_ARM7
	
	define_proc {
	    puts $::cdl_header "#define HAL_PLATFORM_CPU    \"ARM 7TDMI\""
	}
    }

    cdl_component CYGPKG_HAL_ARM_INTEGRATOR_ARM9 {
	display "ARM 9 specialization"
	active_if  CYGPKG_HAL_ARM_ARM9
	calculated CYGPKG_HAL_ARM_ARM9
	
	requires    CYGPKG_HAL_ARM_ARM9_ARM966E
	
	define_proc {
	    puts $::cdl_header "#define HAL_PLATFORM_CPU    \"ARM 9\""
	}
	
    }
    
    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        legal_values  {"RAM" "ROM" "ROMRAM"}
        default_value {"RAM"}
	no_define
	define -file system.h CYG_HAL_STARTUP
        description   "
            When targetting the INTEGRATOR eval board it is possible to build
            the system for either RAM bootstrap or ROM bootstrap(s). Select
            'ram' when building programs to load into RAM using onboard
            debug software such as Angel or eCos GDB stubs.  Select 'rom'
            when building a stand-alone application which will be put
            into ROM."

    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_DEFAULT {
        display      "Default console channel."
        flavor       data
        calculated   0
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD {
        display       "Diagnostic serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 115200
        default_value 38400
        description   "
            This option selects the baud rate used for the diagnostic port.
            Note: this should match the value chosen for the GDB port if the
            diagnostic and GDB port are the same."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_BAUD {
        display       "GDB serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 115200
        default_value 38400
        description   "
            This option controls the baud rate used for the GDB connection."
    }

    cdl_option CYGHWR_HAL_ARM_INTEGRATOR_DIAG_LEDS {
        display          "Enable use of PPx LEDs"
        default_value    1
        description      "
            Enabling this option causes eCos to flash the LEDs during
            early board initialization. See vectors.S for
            details. Before calling cyg_start, PP0 is switched on,
            PP1-3 are switched off. The application code can use the
            function hal_diag_led() to control the LEDs after this
            point."
   }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
        display      "Number of communication channels on the board"
        flavor       data
        calculated   2
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
        display          "Debug serial port"
        active_if        CYGPRI_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_CONFIGURABLE
        flavor 		 data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
            The INTEGRATOR board has two serial ports. This option
            chooses which port will be used to connect to a host
            running GDB."
     }

     cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
         display          "Diagnostic serial port"
         active_if        CYGPRI_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_CONFIGURABLE
         flavor data
         legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
         default_value    CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_DEFAULT
         description      "
            The INTEGRATOR board has two serial ports.  This option
            chooses which port will be used for diagnostic output."
     }

    # Real-time clock/counter specifics
    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants"
        flavor        none
    
        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            calculated    1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            calculated    100
        }
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
           calculated    12500
        }
    }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        parent  CYGPKG_NONE
        description   "
	    Global build options including control over
	    compiler flags, linker flags and choice of toolchain."


        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { CYGHWR_THUMB ? "thumb-elf" : "arm-elf" }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { 
		CYGPKG_HAL_ARM_INTEGRATOR_ARM9 ? "-mcpu=arm9 -Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority" :
		 "-mcpu=arm7tdmi -Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -g -O2 -fno-schedule-insns -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority"
	     }
		 
            description   "
                This option controls the global compiler flags which are used to
                compile all packages by default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value {
		CYGPKG_HAL_ARM_INTEGRATOR_ARM9 ? "-Wl,-Map,map -mcpu=arm9 -g -nostdlib -Wl,--gc-sections -Wl,-static" :
		"-Wl,-Map,map -mcpu=arm7tdmi -g -nostdlib -Wl,--gc-sections -Wl,-static" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }

        cdl_option CYGBLD_BUILD_GDB_STUBS {
            display "Build GDB stub ROM image"
            default_value 0
            requires CYGBLD_BUILD_COMMON_GDB_STUBS
            requires { CYG_HAL_STARTUP != "RAM" }
            requires CYGSEM_HAL_ROM_MONITOR
            requires CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT
            requires CYGDBG_HAL_DEBUG_GDB_THREAD_SUPPORT
            requires ! CYGDBG_HAL_COMMON_INTERRUPTS_SAVE_MINIMUM_CONTEXT
            requires ! CYGDBG_HAL_COMMON_CONTEXT_SAVE_MINIMUM
            no_define
            description "
                This option enables the building of the GDB stubs for the
                board. The address of the ELF headers in the image are
                adjusted to ensure loading at an address in memory used
                by the flash tool."

            make -priority 320 {
                <PREFIX>/bin/gdb_module.bin : <PREFIX>/bin/gdb_module.img
                @mv $< $(<:.img=.elf)
                $(OBJCOPY) --strip-debug --change-addresses=0xFC060000 $(<:.img=.elf) $<
                $(OBJCOPY) -O binary $(<:.img=.elf) $@
            }
        }

        cdl_option CYGBLD_BUILD_FLASH_TOOL {
            display "Build flash programming tool"
            default_value 0
            requires { CYG_HAL_STARTUP == "RAM" }
            requires CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL == 1
            requires CYGPKG_LIBC
            requires CYGPKG_KERNEL
            no_define
            description "This option enables the building of the flash programming tool for copying the GDB stubs into flash memory."
            make -priority 320 {
                <PREFIX>/bin/prog_flash.img : <PACKAGE>/src/prog_flash.c
                @sh -c "mkdir -p src $(dir $@)"
                $(CC) -c $(INCLUDE_PATH) -Wp,-MD,deps.tmp -I$(dir $<) $(CFLAGS) -o src/prog_flash.o $<
                @echo $@ ": \\" > $(notdir $@).deps
                @echo $(wildcard $(PREFIX)/lib/*) " \\" >> $(notdir $@).deps
                @tail +2 deps.tmp >> $(notdir $@).deps
                @echo >> $(notdir $@).deps
                @rm deps.tmp
                $(CC) $(LDFLAGS) -L$(PREFIX)/lib -Ttarget.ld -o $@ src/prog_flash.o
            }
        }

        cdl_option CYGBLD_BUILD_FLASH_TOOL_BE {
            display "Build flash programming tool for BE images on LE boards"
            default_value 0
            requires { CYG_HAL_STARTUP == "RAM" }
            requires CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL == 1
            requires CYGPKG_LIBC
            requires CYGPKG_KERNEL
            no_define
            description "This option enables the building of the flash
                         programming tool for copying the GDB stubs
                         into flash memory. The tool built by enabling
                         this option must be used when programming BE
                         images on LE boards."
            make -priority 320 {
                <PREFIX>/bin/prog_flash_BE_image_LE_system.img : <PACKAGE>/src/prog_flash.c
                @sh -c "mkdir -p src $(dir $@)"
                $(CC) -DBE_IMAGE -c $(INCLUDE_PATH) -Wp,-MD,deps.tmp -I$(dir $<) $(CFLAGS) -o src/prog_flash_be.o $<
                @echo $@ ": \\" > $(notdir $@).deps
                @echo $(wildcard $(PREFIX)/lib/*) " \\" >> $(notdir $@).deps
                @tail +2 deps.tmp >> $(notdir $@).deps
                @echo >> $(notdir $@).deps
                @rm deps.tmp
                $(CC) $(LDFLAGS) -L$(PREFIX)/lib -Ttarget.ld -o $@ src/prog_flash_be.o
            }
        }
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { CYG_HAL_STARTUP == "RAM"    ? "arm_integrator_ram" : \
		     CYG_HAL_STARTUP == "ROMRAM" ? "arm_integrator_romram" : \
                                                   "arm_integrator_rom" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { CYG_HAL_STARTUP == "RAM"    ? "<pkgconf/mlt_arm_integrator_ram.ldi>" : \
			 CYG_HAL_STARTUP == "ROMRAM" ? "<pkgconf/mlt_arm_integrator_romram.ldi>" : \
                                                       "<pkgconf/mlt_arm_integrator_rom.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { CYG_HAL_STARTUP == "RAM"    ? "<pkgconf/mlt_arm_integrator_ram.h>" : \
			 CYG_HAL_STARTUP == "ROMRAM" ? "<pkgconf/mlt_arm_integrator_romram.h>" : \
                                                       "<pkgconf/mlt_arm_integrator_rom.h>" }
        }
    }


    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP != "RAM" }
        description   "
            Enable this option if this program is to be used as a ROM monitor,
            i.e. applications will be loaded into RAM on the board, and this
            ROM monitor may process exceptions or interrupts generated from the
            application. This enables features such as utilizing a separate
            interrupt stack when exceptions are generated."
    }

    cdl_component CYGPKG_CYGMON_HAL_OPTIONS {
        display       "CygMon HAL options"
        flavor        none
        no_define
        parent        CYGPKG_CYGMON
        active_if     CYGPKG_CYGMON
        description   "
            This option also lists the target's requirements for a valid CygMon
            configuration."

        cdl_option CYGBLD_BUILD_CYGMON_BIN {
            display       "Build CygMon ROM binary image"
            active_if     CYGBLD_BUILD_CYGMON
            default_value 1
            no_define
            description "This option enables the conversion of the CygMon ELF
                         image to a binary image suitable for ROM programming."
    
            make -priority 325 {
                <PREFIX>/bin/cygmon.bin : <PREFIX>/bin/cygmon.elf
                $(OBJCOPY) --strip-debug --change-addresses=0xFC060000 $< $(@:.bin=.img) 
                $(OBJCOPY) -O srec $< $(@:.bin=.srec)
                $(OBJCOPY) -O binary $< $@
            }
        }
    }

    cdl_option CYGSEM_HAL_USE_ROM_MONITOR {
         display       "Work with a ROM monitor"
         flavor        booldata
         legal_values  { "Generic" "GDB_stubs" }
         default_value { CYG_HAL_STARTUP == "RAM" ? "GDB_stubs" : 0 }
         parent        CYGPKG_HAL_ROM_MONITOR
         requires      { CYG_HAL_STARTUP == "RAM" }
         description   "
             Support can be enabled for different varieties of ROM monitor.
             This support changes various eCos semantics such as the encoding
             of diagnostic output, or the overriding of hardware interrupt
             vectors.
             Firstly there is \"Generic\" support which prevents the HAL
             from overriding the hardware vectors that it does not use, to
             instead allow an installed ROM monitor to handle them. This is
             the most basic support which is likely to be common to most
             implementations of ROM monitor.
             \"GDB_stubs\" provides support when GDB stubs are included in
             the ROM monitor or boot ROM."
     }

    cdl_component CYGPKG_REDBOOT_HAL_OPTIONS {
        display       "Redboot HAL options"
        flavor        none
        no_define
        parent        CYGPKG_REDBOOT
        active_if     CYGPKG_REDBOOT
        description   "
            This option lists the target's requirements for a valid Redboot
            configuration."
    
	requires      { !CYGPKG_REDBOOT_FLASH || (CYGBLD_REDBOOT_MIN_IMAGE_SIZE == 0x40000) }
	requires      { !CYGOPT_REDBOOT_FIS_REDBOOT_BACKUP }

        cdl_option CYGBLD_BUILD_REDBOOT_BIN_ROM {
            display       "Build Redboot ROM startup ROM binary image"
            active_if     { CYGBLD_BUILD_REDBOOT && CYG_HAL_STARTUP == "ROM" }
            default_value 1
            no_define
            description "This option enables the conversion of the Redboot ELF
                         image to S-Record and binary image suitable for ROM
                         programming."
    
            make -priority 325 {
                <PREFIX>/bin/redboot.bin : <PREFIX>/bin/redboot.elf
                $(OBJCOPY) --strip-debug $< $(@:.bin=.img) 
                $(OBJCOPY) -O srec --gap-fill 0 $< $(@:.bin=.srec)
                $(OBJCOPY) -O binary $< $@
            }
        }

        cdl_option CYGBLD_BUILD_REDBOOT_BIN_ROMRAM {
            display       "Build Redboot ROMRAM startup ROM binary image"
            active_if     { CYGBLD_BUILD_REDBOOT && CYG_HAL_STARTUP == "ROMRAM" }
            default_value 1
            no_define
            description "This option enables the conversion of the Redboot ELF
                         image to S-Record and binary images suitable for ROM
                         programming."
    
            make -priority 325 {
                <PREFIX>/bin/redboot.bin : <PREFIX>/bin/redboot.elf
                $(OBJCOPY) --strip-debug $< $(@:.bin=.img) 
                $(OBJCOPY) -O srec --adjust-vma 0x24000000 --gap-fill 0 $< $(@:.bin=.srec)
                $(OBJCOPY) -O binary $< $@
            }
        }


    }
}
