# ====================================================================
#
#      edb7xxx_eth_drivers.cdl
#
#      Ethernet drivers - platform dependent support for Cirrus Logic
#                         EDB7xxx family of development boards
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Original data:  gthomas
# Contributors:
# Date:           2000-01-25
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_ARM_EDB7XXX {
    display       "Cirrus Logic ethernet driver for EP7xxx boards"

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_HAL_ARM_EDB7XXX

    implements    CYGHWR_NET_DRIVERS
    implements    CYGHWR_NET_DRIVER_ETH0
    include_dir   .
    include_files ; # none _exported_ whatsoever
    description   "Ethernet driver for Cirrus Logic EP7xxx based
                  development boards."
    compile       -library=libextras.a if_edb7xxx.c

    cdl_component CYGSEM_ARM_EDB7XXX_SET_ESA {
        display       "Set the ethernet station address"
        flavor        bool
        default_value 0
        description   "Enabling this option will allow the ethernet
          station address to be forced to the value set by the
          configuration.  This may be required if the hardware does
          not include a serial EEPROM for the ESA."

        cdl_option CYGDAT_ARM_EDB7XXX_ESA {
          display       "The ethernet station address"
          flavor        data
          default_value {"{0x08, 0x88, 0x12, 0x34, 0x56, 0x78}"}
          description   "The ethernet station address"
        }
    }

    cdl_component CYGPKG_DEVS_ETH_ARM_EDB7XXX_OPTIONS {
        display "Cirrus Logic ethernet driver build options"
        flavor  none
	no_define

        cdl_option CYGPKG_DEVS_ETH_ARM_EDB7XXX_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building the Cirrus Logic ethernet driver package.
                These flags are used in addition
                to the set of global flags."
        }
    }
}

