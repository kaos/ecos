# ====================================================================
#
#      io_flash.cdl
#
#      eCos IO configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Original data:  gthomas
# Contributors:
# Date:           2000-07-06
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_IO_FLASH {
    display       "FLASH device drivers"
    include_dir   cyg/io
    description   "
        This option enables drivers for basic I/O services on
        flash devices."
    doc           redirect/ecos-device-drivers.html

    compile       flash.c
 
    define_proc {
	puts $::cdl_header "#include <pkgconf/system.h>"
	puts $::cdl_header "#ifdef CYGDAT_IO_FLASH_DEVICE_HEADER"
	puts $::cdl_header "# include CYGDAT_IO_FLASH_DEVICE_HEADER"
	puts $::cdl_header "#endif "
    }

    cdl_interface CYGHWR_IO_FLASH_DEVICE {
        display       "Hardware FLASH device drivers"
        description   "
            This option enables the hardware device drivers
	    for the current platform."
    }

    cdl_interface CYGHWR_IO_FLASH_BLOCK_LOCKING {
        display       "Hardware can support block locking"
        description   "
            This option will be enabled by devices which can support
            locking (write-protection) of individual blocks."
    }
}
