# ====================================================================
#
#      io_serial.cdl
#
#      eCos IO configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  gthomas
# Contributors:
# Date:           1999-07-07
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_IO_SERIAL {
    display       "Serial device drivers"
    requires      CYGPKG_ERROR
    include_dir   cyg/io
    description   "
        This option enables drivers for basic I/O services on
        serial devices."
    doc           redirect/ecos-device-drivers.html

    compile       -library=libextras.a common/serial.c common/tty.c \
                  common/haldiag.c
    

    cdl_component CYGPKG_IO_SERIAL_TTY {
        display       "TTY-mode serial device drivers"
        flavor        bool
        default_value 1
        description   "
            This option enables the terminal-like device driver 
            used for serial devices that interact with humans,
            such as a system console."
        
        script        tty.cdl
    }

    # -------------------------------------------------------------------------
    cdl_component CYGPKG_IO_SERIAL_ARM_PID {
        display       "ARM PID serial device drivers"
        flavor        bool
        active_if     CYGPKG_HAL_ARM_PID
        default_value 0
        description   "
            This option enables the serial device drivers for the ARM PID."

        compile       -library=libextras.a arm/pid_serial_with_ints.c

        script        ser_arm_pid.cdl
    }

    # -------------------------------------------------------------------------
    cdl_component CYGPKG_IO_SERIAL_ARM_AEB {
        display       "ARM AEB-1 serial device drivers"
        flavor        bool
        active_if     CYGPKG_HAL_ARM_AEB
        default_value 0
        description   "
            This option enables the serial device drivers for the ARM AEB-1."

        compile       -library=libextras.a arm/aeb_serial.c

        script        ser_arm_aeb.cdl
    }

    # -------------------------------------------------------------------------
    cdl_component CYGPKG_IO_SERIAL_ARM_EDB7XXX {
        display       "ARM EDB7XXX serial device drivers"
        flavor        bool
        active_if     CYGPKG_HAL_ARM_EDB7XXX
        default_value 0
        description   "
            This option enables the serial device drivers for the 
	Cirrus Logic EDB7XXX."

        compile       -library=libextras.a arm/edb7xxx_serial.c

        script        ser_arm_edb7xxx.cdl
    }

    # -------------------------------------------------------------------------
    cdl_component CYGPKG_IO_SERIAL_ARM_CMA230 {
        display       "Cogent ARM/CMA230 serial device drivers"
        flavor        bool
        default_value 0
        active_if     CYGPKG_HAL_ARM_CMA230
        description   "
            This option enables the serial device drivers for the Cogent 
            ARM/CMA230."

        compile       -library=libextras.a arm/cma230_serial.c

        script        ser_arm_cma230.cdl
    }

    # -------------------------------------------------------------------------
    cdl_component CYGPKG_IO_SERIAL_POWERPC_COGENT {
        display       "Cogent PowerPC serial device drivers"
        flavor        bool
        active_if     CYGPKG_HAL_POWERPC_COGENT
        default_value 0
        description   "
            This option enables the serial device drivers for the 
            Cogent PowerPC."

        compile       -library=libextras.a powerpc/cogent_serial_with_ints.c

        script        ser_powerpc_cogent.cdl
    }

    # -------------------------------------------------------------------------
    cdl_component CYGPKG_IO_SERIAL_POWERPC_QUICC_SMC {
        display       "PowerPC QUICC/SMC serial device drivers"
        flavor        bool
        active_if     CYGPKG_HAL_QUICC
        default_value 0
        description   "
            This option enables the serial device drivers for the PowerPC 
            QUICC/SMC."

        compile       -library=libextras.a powerpc/quicc_smc_serial.c

        script        ser_quicc_smc.cdl
    }

    # -------------------------------------------------------------------------
    cdl_component CYGPKG_IO_SERIAL_SPARCLITE_SLEB {
        display       "SPARClite SLEB serial device drivers"
        flavor        bool
        active_if     CYGPKG_HAL_SPARCLITE_SLEB
        default_value 0
        description   "
            This option enables the serial device drivers for the 
            SPARClite SLEB."

        compile       -library=libextras.a sparclite/sleb_sdtr.c

        script        ser_sparclite_sleb.cdl
    }

    # -------------------------------------------------------------------------
    cdl_component CYGPKG_IO_SERIAL_TX39_JMR3904 {
        display       "TX39 JMR3904 serial device drivers"
        flavor        bool
        active_if     CYGPKG_HAL_MIPS_TX39_JMR3904
        default_value 0
        description   "
            This option enables the serial device drivers for the TX39 
            JMR3904."

        compile       -library=libextras.a mips/tx3904_serial.c

        script        ser_mips_jmr3904.cdl
    }

    # -------------------------------------------------------------------------
    cdl_component CYGPKG_IO_SERIAL_MIPS_VRC4373 {
        display       "VRC4373 serial device drivers"
        flavor        bool
        active_if     CYGPKG_HAL_MIPS_VR4300_VRC4373
        default_value 0
        description   "
            This option enables the serial device drivers for the VRC4373."

        compile       -library=libextras.a mips/vrc4373_serial.c

        script        ser_mips_vrc4373.cdl
    }

    # -------------------------------------------------------------------------
    # Note: this is not currently tied to a specific board since the
    # ports are "on chip"
    cdl_component CYGPKG_IO_SERIAL_MN10300 {
        display       "MN10300 serial device drivers"
        flavor        bool
        active_if     CYGPKG_HAL_MN10300
        default_value 0
        description   "
            This option enables the serial device drivers for the MN10300."

        compile       -library=libextras.a mn10300/mn10300_serial.c

        script        ser_mn10300.cdl
    }

    # -------------------------------------------------------------------------
    cdl_component CYGPKG_IO_SERIAL_I386_PC {
        display       "PC serial device drivers"
        flavor        bool
        active_if     CYGPKG_HAL_I386_PC
        default_value 0
        description   "
            This option enables the serial device drivers for the PC."

        compile       -library=libextras.a i386/pc_serial.c

        script        ser_i386_pc.cdl
    }

    # -------------------------------------------------------------------------
    cdl_component CYGPKG_IO_SERIAL_SH_EDK7708 {
        display       "SH3 EDK7708 serial device drivers"
        flavor        bool
        active_if CYGPKG_HAL_SH_EDK7708
        default_value 0
        description   "
            This option enables the serial device driver for the Hitachi
            SH3 EDK7708 board."

        compile       -library=libextras.a sh/sh_sci_serial.c

        script        ser_sh_edk7708.cdl
    }

    cdl_component CYGPKG_IO_SERIAL_OPTIONS {
        display "Serial device driver build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_IO_SERIAL_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the serial device drivers. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_IO_SERIAL_CFLAGS_REMOVE {
            display "Supressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the serial device drivers. These flags are removed from
                the set of global flags if present."
        }

        cdl_option CYGPKG_IO_SERIAL_TESTS {
            display "Serial device driver tests"
            flavor  data
            no_define
            calculated { "tests/serial1 tests/serial2 tests/serial3 tests/serial4 tests/serial5 tests/tty1 tests/tty2" }
            description   "
                This option specifies the set of tests for the serial device drivers."
        }
    }
}
