#====================================================================
#
#      ftpclient.cdl
#
#      SNMP library configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      andrew.lunn@ascom.ch
# Original data:  andrew.lunn@ascom.ch
# Contributors:   
# Date:           2001-11-04
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_NET_FTPCLIENT {
    display       "FTP client"
    parent        CYGPKG_NET
    requires      CYGPKG_IO
    requires      { 0 != CYGINT_ISO_STRING_STRFUNCS }
    requires      { 0 != CYGINT_ISO_STRING_MEMFUNCS }
    requires      { 0 != CYGINT_ISO_STDLIB_STRCONV }
    requires      { 0 != CYGINT_ISO_STDIO_FORMATTED_IO }
    requires      { 0 != CYGINT_ISO_STRING_STRFUNCS }
    requires      { 0 != CYGINT_ISO_ERRNO }
    requires      { 0 != CYGINT_ISO_ERRNO_CODES }
    requires      { 0 != CYGINT_ISO_CTYPE }
    requires      CYGPKG_NET
    description   "
        FTP client support. Provides ftp_put and ftp_get to put a file
        onto a remote FTP server and get a file from a remote server. 
        Only binary more is supported."

    compile       ftpclient.c

    cdl_component CYGPKG_NET_FTPCLIENT_OPTIONS {
        display "FTP client build options"
        flavor  none
	no_define

        cdl_option CYGPKG_NET_FTPCLIENT_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building the FTP client package. These flags are used 
                in addition to the set of global flags."
        }

        cdl_option CYGPKG_NET_FTPCLIENT_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the FTP client package. These flags are removed from
                the set of global flags if present."
        }
    }
    cdl_option CYGPKG_NET_FTPCLIENT_TESTS {
        display "FTP Client tests"
        flavor  data
        no_define
        calculated { "tests/ftpclient1.c"}
            description   "
                This option specifies the set of tests for the ftpclient package."
    }
}

