# ====================================================================
#
#      atlas_eth_drivers.cdl
#
#      Ethernet drivers - platform dependent support for MIPS Atlas
#                         board using a Philips SAA9730 IO chip.
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
# -------------------------------------------
# This file is part of eCos, the Embedded Configurable Operating System.
# Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
#
# eCos is free software; you can redistribute it and/or modify it under
# the terms of the GNU General Public License as published by the Free
# Software Foundation; either version 2 or (at your option) any later version.
#
# eCos is distributed in the hope that it will be useful, but WITHOUT ANY
# WARRANTY; without even the implied warranty of MERCHANTABILITY or
# FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
# for more details.
#
# You should have received a copy of the GNU General Public License along
# with eCos; if not, write to the Free Software Foundation, Inc.,
# 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
#
# As a special exception, if other files instantiate templates or use macros
# or inline functions from this file, or you compile this file and link it
# with other works to produce a work based on this file, this file does not
# by itself cause the resulting work to be covered by the GNU General Public
# License. However the source code for this file must still be made available
# in accordance with section (3) of the GNU General Public License.
#
# This exception does not invalidate any other reasons why a work based on
# this file might be covered by the GNU General Public License.
#
# Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
# at http://sources.redhat.com/ecos/ecos-license
# -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      msalter
# Original data:  msalter
# Contributors:
# Date:           2000-12-04
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_MIPS_ATLAS {
    display       "MIPS Atlas ethernet driver"

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_HAL_MIPS_ATLAS

    implements    CYGHWR_NET_DRIVERS
    implements    CYGHWR_NET_DRIVER_ETH0
    include_dir   .
    include_files ; # none _exported_ whatsoever
    description   "Ethernet driver for MIPS Atlas boards w/ SAA9730."
    compile       -library=libextras.a if_atlas.c if_buffers.S

    cdl_component CYGSEM_MIPS_ATLAS_SET_ESA {
        display       "Set the ethernet station address"
        flavor        bool
        default_value 0
        description   "Enabling this option will allow the ethernet
          station address to be forced to the value set by the
          configuration.  This may be required if the hardware does
          not include a serial EEPROM for the ESA."

        cdl_option CYGDAT_MIPS_ATLAS_ESA {
          display       "The ethernet station address"
          flavor        data
          default_value {"{0x00, 0xd0, 0xa0, 0x00, 0x00, 0x10}"}
          description   "The ethernet station address"
        }
    }

    cdl_component CYGPKG_DEVS_ETH_MIPS_ATLAS_OPTIONS {
        display "MIPS Atlas ethernet driver build options"
        flavor  none
	no_define

        cdl_option CYGPKG_DEVS_ETH_ARM_ATLAS_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building the MIPS Atlas ethernet driver package.
                These flags are used in addition
                to the set of global flags."
        }
    }
}

