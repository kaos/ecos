# ====================================================================
#
#      eth_drivers.cdl
#
#      Ethernet drivers - platform independent support
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Original data:  gthomas
# Contributors:
# Date:           2000-01-25
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_IO_ETH_DRIVERS {
    display       "Common ethernet support"
    include_dir   .
    parent        CYGPKG_IO
    description   "Platform independent ethernet drivers"

    cdl_component CYGPKG_IO_ETH_DRIVERS_NET {
        display       "Support for standard eCos TCP/IP stack."
        flavor        bool
        active_if     CYGPKG_NET
        no_define
        default_value 1
        compile       net/eth_drv.c
    }

    cdl_component CYGPKG_IO_ETH_DRIVERS_STAND_ALONE {
        display       "Support for stand-alone network stack."
        flavor        bool
        active_if     !CYGPKG_NET
        default_value 1
        no_define
        compile       stand_alone/eth_drv.c

        cdl_option CYGNUM_IO_ETH_DRIVERS_NUM_PKT {
            display          "Number of \[network\] buffers"
            flavor           data
            default_value    16
            legal_values     2 to 32
            description      "
               This option is used to allocate space to buffer incoming network
               packets.  These buffers are used to hold data until they can be
               logically processed by higher layers."
        }

        cdl_option CYGSEM_IO_ETH_DRIVERS_WARN {
            display          "Show driver warnings"
            flavor           bool
            default_value    0
            description      "
               Selecting this option will allows the stand-alone ethernet driver
               to display warnings on the system console when incoming network
               packets are being discarded due to lack of buffer space."
        }

        cdl_option CYGSEM_IO_ETH_DRIVERS_DEBUG {
            display          "Print driver debug information"
            flavor           bool
            default_value    0
            description      "
               Selecting this option will enable the stand-alone driver to print
               lots of information.  Useful only when getting a low-level hardware
               driver to work."
        }
    }

    cdl_component CYGPKG_IO_ETH_DRIVERS_OPTIONS {
        display "Common ethernet support build options"
        flavor  none
	no_define

        cdl_option CYGPKG_IO_ETH_DRIVERS_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building the common ethernet support package. These flags are used in addition
                to the set of global flags."
        }
    }
}
