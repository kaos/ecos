# ====================================================================
#
#      hal_arm_arm9_aaed2000.cdl
#
#      Agilent AAED2000 platform HAL package configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Original data:  gthomas
# Contributors:
# Date:           2001-10-27
#
#####DESCRIPTIONEND####
#
# ====================================================================
cdl_package CYGPKG_HAL_ARM_ARM9_AAED2000 {
    display       "Agilent Aaed2000 evaluation board"
    parent        CYGPKG_HAL_ARM_ARM9
    requires      CYGPKG_HAL_ARM_ARM9_ARM920T
    hardware
    include_dir   cyg/hal
    define_header hal_arm_arm9_aaed2000.h
    description   "
        This HAL platform package provides generic
        support for the Agilent based board, known as 'aaed2000'."

    compile       aaed2000_misc.c hal_diag.c kbd_drvr.c

    implements    CYGINT_HAL_DEBUG_GDB_STUBS
    implements    CYGINT_HAL_DEBUG_GDB_STUBS_BREAK
    implements    CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT
    implements    CYGINT_HAL_PLF_IF_INIT


    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H   <pkgconf/hal_arm.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_VARIANT_H  <pkgconf/hal_arm_arm9.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_arm_arm9_aaed2000.h>"

        puts $::cdl_header "#define HAL_PLATFORM_CPU    \"ARM9\""
        puts $::cdl_header "#define HAL_PLATFORM_BOARD  \"AAED2000 system\""
        puts $::cdl_header "#define HAL_PLATFORM_EXTRA  \"\[\" __Xstr(CYGHWR_REDBOOT_BOOTMONITOR) \"\]\" "
        puts $::cdl_header "#define HAL_PLATFORM_MACHINE_TYPE  106"
    }

    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        default_value {"RAM"}
        legal_values  {"RAM" "ROM" "ROMRAM" }
	no_define
	define -file system.h CYG_HAL_STARTUP
        description   "
           When targetting the Aaed2000 eval board it is possible to build
           the system for either RAM bootstrap or ROM bootstrap(s). Select
           'ram' when building programs to load into RAM using eCos GDB
           stubs.  Select 'rom' when building a stand-alone application
           which will be put into ROM, or for the special case of
           building the eCos GDB stubs themselves."
    }

    cdl_component CYGNUM_HAL_ARM_AAED2000_CLOCK {
        display       "Board (CPU and bus) speed"
        flavor data
        legal_values  {"150/75MHz" "166/83MHz"}
        default_value {"150/75MHz"}
        description   "
            This option controls the CPU and bus frequencies. It
            does so by presetting the PLL details when one of the
            frequency combinations are selected. It's also possible
            to customize the PLL values by selecting 'Custom'
            and adjusting the options accordingly. See the 'Clock and Control'
            section of the CPU manual for further information."

        # Note: there are options for these settings, even though they
        # are compute. That's because I initially thought the cpu/bus
        # speed could be calculated properly - for now they are also
        # just set as a result of the _CLOCK choice.
        # See table 5-7 in the manual for the setting of these parameters.
        cdl_option CYGNUM_HAL_ARM_AAED2000_CLOCK_REF {
            display       "CPU clock reference clock (crystal)"
            flavor        data
            calculated    14745600
            description   "
                This is the CPU reference clock. It is 14.7456MHz and
                cannot be changed."
        }

        cdl_option CYGNUM_HAL_ARM_AAED2000_CLOCK_HCLKDIV {
            display       "CPU clock HCLKDIV"
            flavor        data
            calculated    { CYGNUM_HAL_ARM_AAED2000_CLOCK == "150/75MHz" ? 1 :
                            CYGNUM_HAL_ARM_AAED2000_CLOCK == "166/83MHz" ? 1 :
                             0 }
            description   "
                The HCLKDIV value."
        }

        cdl_option CYGNUM_HAL_ARM_AAED2000_CLOCK_PREDIV {
            display       "CPU clock PREDIV"
            flavor        data
            calculated    { CYGNUM_HAL_ARM_AAED2000_CLOCK == "150/75MHz" ? 12 :
                            CYGNUM_HAL_ARM_AAED2000_CLOCK == "166/83MHz" ? 18 :
                             0 }
            description   "
                The PREDIV value."
        }

        cdl_option CYGNUM_HAL_ARM_AAED2000_CLOCK_MAINDIV1 {
            display       "CPU clock MAINDIV1"
            flavor        data
            calculated    { CYGNUM_HAL_ARM_AAED2000_CLOCK == "150/75MHz" ? 13 :
                            CYGNUM_HAL_ARM_AAED2000_CLOCK == "166/83MHz" ? 13 :
                             0 }
            description   "
                The MAINDIV1 value."
        }

        cdl_option CYGNUM_HAL_ARM_AAED2000_CLOCK_MAINDIV2 {
            display       "CPU clock MAINDIV2"
            flavor        data
            calculated    { CYGNUM_HAL_ARM_AAED2000_CLOCK == "150/75MHz" ? 17 :
                            CYGNUM_HAL_ARM_AAED2000_CLOCK == "166/83MHz" ? 28 :
                             0 }
            description   "
                The MAINDIV2 value."
        }

        cdl_option CYGNUM_HAL_ARM_AAED2000_CLOCK_PCLKDIV {
            display       "CPU clock PCLKDIV"
            flavor        data
            calculated    { CYGNUM_HAL_ARM_AAED2000_CLOCK == "150/75MHz" ? 1 :
                            CYGNUM_HAL_ARM_AAED2000_CLOCK == "166/83MHz" ? 1 :
                             0 }
            description   "
                The PCLKDIV value."
        }

        cdl_option CYGNUM_HAL_ARM_AAED2000_CLOCK_PS {
            display       "CPU clock PS"
            flavor        data
            calculated    { CYGNUM_HAL_ARM_AAED2000_CLOCK == "150/75MHz" ? 1 :
                            CYGNUM_HAL_ARM_AAED2000_CLOCK == "166/83MHz" ? 1 :
                             0 }
            description   "
                The PCLKDIV value."
        }


        cdl_option CYGNUM_HAL_ARM_AAED2000_CPU_CLOCK {
            display       "CPU speed"
            flavor        data
            calculated    { CYGNUM_HAL_ARM_AAED2000_CLOCK == "150/75MHz" ? 150890000 :
                            CYGNUM_HAL_ARM_AAED2000_CLOCK == "166/83MHz" ? 165888000 :
                             0 }
            description   "
            This is the actual CPU operating frequency."
        }

        cdl_option CYGNUM_HAL_ARM_AAED2000_BUS_CLOCK {
            display       "Bus speed"
            flavor        data
            calculated    { CYGNUM_HAL_ARM_AAED2000_CLOCK == "150/75MHz" ?  75445000 :
                            CYGNUM_HAL_ARM_AAED2000_CLOCK == "166/83MHz" ?  82944000 :
                             0 }
            description   "
            This is the actual bus operating frequency."
        }
    }


    # Real-time clock/counter specifics
    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants"
        flavor        none
        no_define
    
        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            default_value 1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            default_value 100
        }
        # The timer used runs at 508kHz
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
            default_value ((508000/CYGNUM_HAL_RTC_DENOMINATOR)-1)
        }
    }

    cdl_component CYGSEM_AAED2000_LCD_SUPPORT {
        display        "Support LCD"
        flavor         bool
        default_value  1
        compile        lcd_support.c
        description    "
          Enabling this option will enable the use the LCD as a 
          simple framebuffer, suitable for use with a windowing
          package."

        cdl_option  CYGSEM_AAED2000_LCD_PORTRAIT_MODE {
            display       "LCD portrait mode"
            flavor        bool
            default_value 0
            description   "
                Setting this option will orient the data on the LCD screen
                in portrait (480x640) mode."
        }

        cdl_component CYGSEM_AAED2000_LCD_COMM {
            display        "Support LCD/keyboard for comminication channel"
            active_if      CYGPKG_REDBOOT
            flavor         bool
            default_value  1
            description    "
              Enabling this option will use the LCD and keyboard for a
              communications channel, suitable for RedBoot, etc."

            cdl_option  CYGOPT_AAED2000_LCD_COMM_LOGO {
                display       "RedHat logo location"
                flavor        booldata
                legal_values  { "TOP" "BOTTOM" }
                default_value { "TOP" }
                description   "
                    Use this option to control where the RedHat logo is placed
                    on the LCD screen."
            }
        }
    }
    

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD {
        display       "Diagnostic serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 57600 115200
        default_value 38400
        description   "
            This option selects the baud rate used for the diagnostic port.
            Note: this should match the value chosen for the GDB port if the
            diagnostic and GDB port are the same."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_BAUD {
        display       "GDB serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 57600 115200
        default_value 38400
        description   "
            This option selects the baud rate used for the diagnostic port.
            Note: this should match the value chosen for the GDB port if the
            diagnostic and GDB port are the same."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
        display      "Number of communication channels on the board"
        flavor       data
        calculated   1+CYGSEM_AAED2000_LCD_COMM
    }
 
    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
        display          "Debug serial port"
        active_if        CYGPRI_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_CONFIGURABLE
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
            The aaed2000 board has two serial ports. This option
            chooses which port will be used to connect to a host
            running GDB."
     }

     cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_DEFAULT {
         display      "Default console channel."
         flavor       data
         legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
         calculated   0
     }
 
     cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
         display          "Diagnostic serial port"
         active_if        CYGPRI_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_CONFIGURABLE
         flavor data
         legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
         default_value    CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_DEFAULT
         description      "
            The aaed2000 board has two serial ports.  This option
            chooses which port will be used for diagnostic output."
     }
 
    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        no_define
        description   "
	    Global build options including control over
	    compiler flags, linker flags and choice of toolchain."


        parent  CYGPKG_NONE

        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "arm-eabi"}
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { "-mcpu=arm9 -Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority" }
            description   "
                This option controls the global compiler flags which are used to
                compile all packages by default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { "-Wl,--gc-sections -Wl,-static -g -O2 -nostdlib" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }

        cdl_option CYGBLD_BUILD_GDB_STUBS {
            display "Build GDB stub ROM image"
            default_value 0
            requires { CYG_HAL_STARTUP == "ROM" }
            requires CYGSEM_HAL_ROM_MONITOR
            requires CYGBLD_BUILD_COMMON_GDB_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT
            requires CYGDBG_HAL_DEBUG_GDB_THREAD_SUPPORT
            requires ! CYGDBG_HAL_COMMON_INTERRUPTS_SAVE_MINIMUM_CONTEXT
            requires ! CYGDBG_HAL_COMMON_CONTEXT_SAVE_MINIMUM
            no_define
            description "
                This option enables the building of the GDB stubs for the
                board. The common HAL controls takes care of most of the
                build process, but the final conversion from ELF image to
                binary data is handled by the platform CDL, allowing
                relocation of the data if necessary."

            make -priority 320 {
                <PREFIX>/bin/gdb_module.srec : <PREFIX>/bin/gdb_module.img
                $(OBJCOPY) --remove-section=.fixed_vectors $< gdb_module.tmp
                $(OBJCOPY) -O srec --change-address 0x10000000 gdb_module.tmp $@
            }
        }
    }

    cdl_component CYGPKG_HAL_ARM_ARM9_AAED2000_OPTIONS {
        display "ARM9/AAED2000 build options"
        flavor  none
        no_define
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_HAL_ARM_ARM9_AAED2000_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the ARM9 AAED2000 HAL. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_HAL_ARM_ARM9_AAED2000_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the ARM9 AAED2000 HAL. These flags are removed from
                the set of global flags if present."
        }

        cdl_option CYGPKG_HAL_ARM_ARM9_AAED2000_TESTS {
            display "ARM9/AAED2000 tests"
            flavor  data
            no_define
            calculated { "" }
            description   "
                This option specifies the set of tests for the ARM9 Aaed2000 HAL."
        }
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { CYG_HAL_STARTUP == "RAM" ? "arm_arm9_aaed2000_ram" : \
	             CYG_HAL_STARTUP == "ROM" ? "arm_arm9_aaed2000_rom" : \
                                                "arm_arm9_aaed2000_romram" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_arm9_aaed2000_ram.ldi>" : \
                         CYG_HAL_STARTUP == "ROM" ? "<pkgconf/mlt_arm_arm9_aaed2000_rom.ldi>" : \
                                                    "<pkgconf/mlt_arm_arm9_aaed2000_romram.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_arm9_aaed2000_ram.h>" : \
                         CYG_HAL_STARTUP == "ROM" ? "<pkgconf/mlt_arm_arm9_aaed2000_rom.h>" : \
                                                    "<pkgconf/mlt_arm_arm9_aaed2000_romram.h>" }
        }
    }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "ROM" || CYG_HAL_STARTUP == "ROMRAM" }
        description   "
            Enable this option if this program is to be used as a ROM monitor,
            i.e. applications will be loaded into RAM on the board, and this
            ROM monitor may process exceptions or interrupts generated from the
            application. This enables features such as utilizing a separate
            interrupt stack when exceptions are generated."
    }

    cdl_option CYGSEM_HAL_USE_ROM_MONITOR {
         display       "Work with a ROM monitor"
         flavor        booldata
         legal_values  { "Generic" "GDB_stubs" }
         default_value { CYG_HAL_STARTUP == "RAM" ? "GDB_stubs" : 0 }
         parent        CYGPKG_HAL_ROM_MONITOR
         requires      { CYG_HAL_STARTUP == "RAM" }
         description   "
             Support can be enabled for different varieties of ROM monitor.
             This support changes various eCos semantics such as the encoding
             of diagnostic output, or the overriding of hardware interrupt
             vectors.
             Firstly there is \"Generic\" support which prevents the HAL
             from overriding the hardware vectors that it does not use, to
             instead allow an installed ROM monitor to handle them. This is
             the most basic support which is likely to be common to most
             implementations of ROM monitor.
             \"GDB_stubs\" provides support when GDB stubs are included in
             the ROM monitor or boot ROM."
     }

    cdl_component CYGPKG_REDBOOT_HAL_OPTIONS {
        display       "Redboot HAL options"
        flavor        none
        no_define
        parent        CYGPKG_REDBOOT
        active_if     CYGPKG_REDBOOT
        description   "
            This option lists the target's requirements for a valid Redboot
            configuration."

        # The backup image is not needed, since ROMRAM is the normal
        # RedBoot startup type.
        requires {!CYGPKG_REDBOOT_FLASH || CYGOPT_REDBOOT_FIS_REDBOOT_BACKUP == 0}

        # RedBoot details
        requires { CYGPKG_REDBOOT_ARM_LINUX_EXEC }
        requires { CYGHWR_REDBOOT_ARM_LINUX_EXEC_ADDRESS_DEFAULT == 0xf0008000 }
        define_proc {
            puts $::cdl_header "#define CYGHWR_REDBOOT_ARM_TRAMPOLINE_ADDRESS 0x00001f00"
        }

        cdl_option CYGHWR_REDBOOT_BOOTMONITOR {
            display       "Controls where RedBoot is in the boot chain"
            default_value {"Primary"}
            legal_values  {"Primary"}
            flavor        data
            active_if     CYGPKG_REDBOOT_FLASH
            description   "
                This option selects whether RedBoot sits in the boot chain.
                Presently it's only supported as the primary booter."

        }
        cdl_option CYGBLD_BUILD_REDBOOT_BIN {
            display       "Build Redboot ROM binary image"
            active_if     CYGBLD_BUILD_REDBOOT
            default_value 1
            no_define
            description "This option enables the conversion of the Redboot ELF
                         image to the various relocated SREC images needed
                         for flash updating."

            make -priority 325 {
                <PREFIX>/bin/redboot.bin : <PREFIX>/bin/redboot.elf
                $(OBJCOPY) --strip-debug $< $(@:.bin=.img) 
                $(OBJCOPY) -O srec $< $(@:.bin=.srec)
                $(OBJCOPY) -O binary $< $@
            }
        }
    }

}
