# ====================================================================
#
#      spi_lpc2xxx.cdl
#
#      SPI driver for LPC2xxx
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Hans Rosenfeld <rosenfeld@grumpf.hope-2000.org>
# Contributors:   
# Date:           2007-07-12
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_SPI_ARM_LPC2XXX {
    display     "LPC2xxx SPI driver"
    requires    CYGPKG_HAL_ARM_LPC2XXX

    parent      CYGPKG_IO_SPI
    active_if   CYGPKG_IO_SPI

    include_dir cyg/io
    compile     spi_lpc2xxx.cxx

    cdl_option CYGPKG_DEVS_SPI_ARM_LPC2XXX_BUS0 {
        display       "Enable SPI interface 0"
        flavor        bool
        default_value 1
        description   "The LPC2xxx controllers contain two SPI interfaces.
                       Enable this option to get support for SPI interface 0."
    }

    cdl_option CYGPKG_DEVS_SPI_ARM_LPC2XXX_BUS1 {
        display       "Enable SPI interface 1"
        flavor        bool
        default_value 1
        description   "The LPC2xxx controllers contain two SPI interfaces.
                       Enable this option to get support for SPI interface 1."
    }
}
