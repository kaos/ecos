#====================================================================
#
#      ftpclient.cdl
#
#      SNMP library configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
# -------------------------------------------
# This file is part of eCos, the Embedded Configurable Operating System.
# Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
#
# eCos is free software; you can redistribute it and/or modify it under
# the terms of the GNU General Public License as published by the Free
# Software Foundation; either version 2 or (at your option) any later version.
#
# eCos is distributed in the hope that it will be useful, but WITHOUT ANY
# WARRANTY; without even the implied warranty of MERCHANTABILITY or
# FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
# for more details.
#
# You should have received a copy of the GNU General Public License along
# with eCos; if not, write to the Free Software Foundation, Inc.,
# 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
#
# As a special exception, if other files instantiate templates or use macros
# or inline functions from this file, or you compile this file and link it
# with other works to produce a work based on this file, this file does not
# by itself cause the resulting work to be covered by the GNU General Public
# License. However the source code for this file must still be made available
# in accordance with section (3) of the GNU General Public License.
#
# This exception does not invalidate any other reasons why a work based on
# this file might be covered by the GNU General Public License.
#
# Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
# at http://sources.redhat.com/ecos/ecos-license
# -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      andrew.lunn@ascom.ch
# Original data:  andrew.lunn@ascom.ch
# Contributors:   
# Date:           2001-11-04
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_NET_FTPCLIENT {
    display       "FTP client"
    parent        CYGPKG_NET
    requires      CYGPKG_IO
    requires      { 0 != CYGINT_ISO_STRING_STRFUNCS }
    requires      { 0 != CYGINT_ISO_STRING_MEMFUNCS }
    requires      { 0 != CYGINT_ISO_STDLIB_STRCONV }
    requires      { 0 != CYGINT_ISO_STDIO_FORMATTED_IO }
    requires      { 0 != CYGINT_ISO_STRING_STRFUNCS }
    requires      { 0 != CYGINT_ISO_ERRNO }
    requires      { 0 != CYGINT_ISO_ERRNO_CODES }
    requires      { 0 != CYGINT_ISO_CTYPE }
    requires      CYGPKG_NET
    description   "
        FTP client support. Provides ftp_put and ftp_get to put a file
        onto a remote FTP server and get a file from a remote server. 
        Only binary more is supported."

    compile       ftpclient.c

    cdl_component CYGPKG_NET_FTPCLIENT_OPTIONS {
        display "FTP client build options"
        flavor  none
	no_define

        cdl_option CYGPKG_NET_FTPCLIENT_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building the FTP client package. These flags are used 
                in addition to the set of global flags."
        }

        cdl_option CYGPKG_NET_FTPCLIENT_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the FTP client package. These flags are removed from
                the set of global flags if present."
        }
    }
    cdl_option CYGPKG_NET_FTPCLIENT_TESTS {
        display "FTP Client tests"
        flavor  data
        no_define
        calculated { "tests/ftpclient1.c"}
            description   "
                This option specifies the set of tests for the ftpclient package."
    }
}

