# ====================================================================
#
#      hal_arm_cma230.cdl
#
#      Cogent CMA230 board HAL package configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  gthomas
# Contributors:
# Date:           1999-07-01
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_ARM_CMA230 {
    display       "Cogent Computer Systems CMA2xx boards"
    parent        CYGPKG_HAL_ARM
    hardware
    include_dir   cyg/hal
    define_header hal_arm_cma230.h
    description   "
        The cma230 HAL package provides the support needed to run
        eCos on Cogent Computer Systems CMA2xx (CMA230, CMA222) boards."

    compile       hal_diag.c plf_stub.c cma230_misc.c

    implements    CYGINT_HAL_DEBUG_GDB_STUBS
    implements    CYGINT_HAL_DEBUG_GDB_STUBS_BREAK

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H   <pkgconf/hal_arm.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_arm_cma230.h>"
    }

    cdl_option CYGHWR_HAL_ARM_CMA2XX_VARIANT {
        display       "Cogent CMA2xxx processor variant"
        flavor        data
        legal_values  { "CMA230" "CMA222" }
        default_value { "CMA230" }
        description   "
            The processor variant used by the Cogent board."
    }

    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        legal_values  {"RAM" "ROM"}
        default_value {"RAM"}
	no_define
	define -file system.h CYG_HAL_STARTUP
        description   "
            When targetting the CMA230 board it is possible to build
            the system for either RAM bootstrap or ROM bootstrap(s). Select
            'ram' when building programs to load into RAM using onboard
            debug software such as Angel or eCos GDB stubs.  Select 'rom'
            when building a stand-alone application which will be put
            into ROM."
    }

    cdl_option CYGHWR_HAL_ARM_CMA230_DIAG_PORT {
        display       "Diagnostic serial port"
        flavor        data
        legal_values  0 1
        default_value 0
        description   "
            The CMA230 board has two separate serial ports.  This option
            chooses which of these ports will be used."
    }
    
    cdl_option CYGHWR_HAL_ARM_CMA230_DIAG_BAUD {
        display       "Diagnostic serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 115200
        default_value 38400
        description   "
            This option selects the baud rate used for the diagnostic port.
            Note: this should match the value chosen for the GDB port if the
            diagnostic and GDB port are the same."
    }
    
    cdl_option CYGHWR_HAL_ARM_CMA230_GDB_PORT {
        display       "GDB serial port"
        flavor        data
        legal_values  0 1
        default_value 0
        description   "
            The CMA230 board has two separate serial ports.  This option
            chooses which of these ports will be used to connect to a host
            running GDB."
    }

    cdl_option CYGHWR_HAL_ARM_CMA230_GDB_BAUD {
        display       "GDB serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 115200
        default_value 38400
        description   "
            This option controls the baud rate used for the GDB connection."
    }

    # Real-time clock/counter specifics
    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants"
        flavor        none
    
        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            calculated    1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            calculated    100
        }
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
           calculated    5000                    ;# 2us clock
        }
    }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        parent  CYGPKG_NONE
        description   "
	    Global build options including control over
	    compiler flags, linker flags and choice of toolchain."


        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            if {1} {
                default_value { CYGHWR_THUMB ? "thumb-elf" : "arm-elf" }
            } else {
                default_value { "arm-elf" }
            }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            if {1} {
                default_value { CYGHWR_THUMB ? "-mthumb-interwork -Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority" :
                "-mcpu=arm7tdmi -Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority" }
            } else {
                default_value { "-mcpu=arm7tdmi -Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority" }
            }
            description   "
                This option controls the global compiler flags which are used to
                compile all packages by default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGPKG_HAL_ARM_CMA2XX_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { CYGHWR_HAL_ARM_CMA2XX_VARIANT == "CMA222" ? "-D__CMA222" : "" }
            description   "
                This option modifies the set of compiler flags for
                building the Cogent board HAL. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_HAL_ARM_CMA2XX_CFLAGS_REMOVE {
            display "Supressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the Cogent board HAL. These flags are removed from
                the set of global flags if present."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            if {1} {
                default_value { CYGHWR_THUMB ? "-g -nostdlib -Wl,--gc-sections -Wl,-static -mthumb-interwork" :
                                               "-mcpu=arm7tdmi -g -nostdlib -Wl,--gc-sections -Wl,-static" }
            } else {
                default_value { "-mcpu=arm7tdmi -g -nostdlib -Wl,--gc-sections -Wl,-static" }
            }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }

        cdl_option CYGBLD_BUILD_GDB_STUBS {
            display "Build GDB stub ROM image"
            default_value 0
            requires CYGBLD_BUILD_COMMON_GDB_STUBS
            requires { CYG_HAL_STARTUP == "ROM" }
            requires CYGSEM_HAL_ROM_MONITOR
            requires CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
            requires ! CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT
            requires ! CYGDBG_HAL_DEBUG_GDB_THREAD_SUPPORT
            requires ! CYGDBG_HAL_COMMON_INTERRUPTS_SAVE_MINIMUM_CONTEXT
            requires ! CYGDBG_HAL_COMMON_CONTEXT_SAVE_MINIMUM
            no_define
            description "
                This option enables the building of the GDB stubs for the
                board."

            make -priority 320 {
                <PREFIX>/bin/gdb_module.bin : <PREFIX>/bin/gdb_module.img
                @mv $< $(<:.img=.elf)
                $(OBJCOPY) --strip-debug --change-addresses=0x10038000 $(<:.img=.elf) $<
                $(OBJCOPY) -O binary $(<:.img=.elf) $@
            }
        }
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { CYGHWR_HAL_ARM_CMA2XX_VARIANT == "CMA230" ? \
                       (CYG_HAL_STARTUP == "RAM" ? "arm_cma230_ram" : \
                                                   "arm_cma230_rom"): \
                       (CYG_HAL_STARTUP == "RAM" ? "arm_cma222_ram" : \
                                                   "arm_cma222_rom") }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { CYGHWR_HAL_ARM_CMA2XX_VARIANT == "CMA230" ? \
                           (CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_cma230_ram.ldi>" : \
                                                       "<pkgconf/mlt_arm_cma230_rom.ldi>") : \
                           (CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_cma222_ram.ldi>" : \
                                                       "<pkgconf/mlt_arm_cma222_rom.ldi>") }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { CYGHWR_HAL_ARM_CMA2XX_VARIANT == "CMA230" ? \
                           (CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_cma230_ram.h>" : \
                                                       "<pkgconf/mlt_arm_cma230_rom.h>") : \
                           (CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_cma222_ram.h>" : \
                                                       "<pkgconf/mlt_arm_cma222_rom.h>") }
        }
    }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "ROM" }
        description   "
            Enable this option if this program is to be used as a ROM monitor,
            i.e. applications will be loaded into RAM on the board, and this
            ROM monitor may process exceptions or interrupts generated from the
            application. This enables features such as utilizing a separate
            interrupt stack when exceptions are generated."
    }
}
