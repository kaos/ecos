# ====================================================================
#
#      hal_arm_iq80310.cdl
#
#      IQ80310 evaluation board HAL package configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      msalter
# Original data:  
# Contributors:
# Date:           2000-10-09
#
#####DESCRIPTIONEND####
#
# ====================================================================
cdl_package CYGPKG_HAL_ARM_IQ80310 {
    display       "Intel IQ80310 XScale evaluation boards"
    parent        CYGPKG_HAL_ARM
    define_header hal_arm_iq80310.h
    include_dir   cyg/hal
    hardware
    description   "
        The IQ80310 HAL package provides the support needed to run
        eCos on an Intel IQ80310 XScale eval board."

    compile hal_diag.c iq80310_misc.c iq80310_pci.c

    implements    CYGINT_HAL_DEBUG_GDB_STUBS
    implements    CYGINT_HAL_DEBUG_GDB_STUBS_BREAK
    implements    CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT
    implements    CYGINT_HAL_ARM_MEM_REAL_REGION_TOP
    implements    CYGINT_HAL_ARM_ARCH_XSCALE

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H   <pkgconf/hal_arm.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_arm_iq80310.h>"
	puts $::cdl_header "#define HAL_PLATFORM_CPU    \"XScale\""
        puts $::cdl_header "#define HAL_PLATFORM_BOARD  \"IQ80310\""
        puts $::cdl_header "#define HAL_PLATFORM_EXTRA  \"\""
        puts $::cdl_header "#define HAL_ARCH_PROGRAM_NEW_STACK iq80310_program_new_stack"
    }

    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        default_value {"RAM"}
        legal_values  {"RAM" "ROM"}
	no_define
	define -file system.h CYG_HAL_STARTUP
        description   "
           When targetting the IQ80310 eval board it is possible to build
           the system for either RAM bootstrap or ROM bootstrap(s). Select
           'ram' when building programs to load into RAM using onboard
           debug software such as Angel or eCos GDB stubs.  Select 'rom'
           when building a stand-alone application which will be put
           into ROM.  Selection of 'stubs' is for the special case of
           building the eCos GDB stubs themselves."
    }

    cdl_option CYGSEM_HAL_ARM_IQ80310_ARMBOOT {
        display       "Coexist with ARM bootloader"
        flavor        bool
        default_value 0
        description   "
            Enable this option if the ARM bootloader is programmed into
            the FLASH boot sector on the board."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_DEFAULT {
        display      "Default console channel."
        flavor       data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        calculated   0
    }
 
    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
        display      "Number of communication channels on the board"
        flavor       data
        calculated   2
    }
 
    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
        display          "Debug serial port"
        active_if        CYGPRI_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_CONFIGURABLE
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
            This option chooses which port will be used to connect to a host
            running GDB."
     }
 
     cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
         display          "Diagnostic serial port"
         active_if        CYGPRI_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_CONFIGURABLE
         flavor data
         legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
         default_value    CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_DEFAULT
         description      "
            The EBSA285 board has only one serial port.  This option
            chooses which port will be used for diagnostic output."
     }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD {
        display       "Diagnostic serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 57600 115200
        default_value 115200
        description   "
            This option selects the baud rate used for the diagnostic port.
            Note: this should match the value chosen for the GDB port if the
            diagnostic and GDB port are the same."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_BAUD {
        display       "GDB serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 57600 115200
        default_value 115200
        description   "
            This option selects the baud rate used for the GDB port."
    }

    # Real-time clock/counter specifics
    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants"
        flavor        none
    
        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            calculated    1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            calculated    100
        }
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
            calculated    330000        ;# External timer is 33MHz
        }
    }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        description   "
	    Global build options including control over
	    compiler flags, linker flags and choice of toolchain."


        parent  CYGPKG_NONE

        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "arm-elf" }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { "-mcpu=xscale -Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority -mapcs-frame" }
            description   "
                This option controls the global compiler flags which are used to
                compile all packages by default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { "-mcpu=xscale -Wl,--gc-sections -Wl,-static -g -O2 -nostdlib" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }

        cdl_option CYGBLD_BUILD_GDB_STUBS {
            display "Build GDB stub ROM image"
            default_value 0
            requires { CYG_HAL_STARTUP == "ROM" }
            requires CYGSEM_HAL_ROM_MONITOR
            requires CYGBLD_BUILD_COMMON_GDB_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT
            requires CYGDBG_HAL_DEBUG_GDB_THREAD_SUPPORT
            requires ! CYGDBG_HAL_COMMON_INTERRUPTS_SAVE_MINIMUM_CONTEXT
            requires ! CYGDBG_HAL_COMMON_CONTEXT_SAVE_MINIMUM
            no_define
            description "
                This option enables the building of the GDB stubs for the
                board. The common HAL controls takes care of most of the
                build process, but the final conversion from ELF image to
                binary data is handled by the platform CDL, allowing
                relocation of the data if necessary."

            make -priority 320 {
                <PREFIX>/bin/gdb_module.bin : <PREFIX>/bin/gdb_module.img
                $(OBJCOPY) -O binary $< $@
            }
        }
    }

    cdl_option CYGNUM_HAL_BREAKPOINT_LIST_SIZE {
        display       "Number of breakpoints supported by the HAL."
        flavor        data
        default_value 32
        description   "
            This option determines the number of breakpoints supported by the HAL."
    }

    cdl_component CYGPKG_HAL_ARM_IQ80310_OPTIONS {
        display "XScale IQ80310 build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."

	cdl_option CYGSEM_HAL_ARM_IQ80310_BTB {
            display       "Enable Branch Target Buffer"
            flavor        bool
            default_value 0
            description   "
                Enable this option to turn on the IQ80200 Branch Target Buffer
                which is used for branch prediction. This is turned off by
                default because of CPU errata which may cause thumb branches
                to execute improperly on A-step CPUs. Normal ARM programs are
                not affected by this errata, so enabling this option for
                ARM-only applications may improve program performance."
        }

	cdl_option CYGSEM_HAL_ARM_IQ80310_CLEAR_PCI_RETRY {
            display       "Have RedBoot clear PCI Retry bit"
            flavor        bool
            default_value 1
            description   "
                This option controls whether or not RedBoot allows the host PC
                to completely boot. In some cases, you may not want to allow
                this if RedBoot is used to automatically launch an application
                which needs to run some setup code before allowing the PC to
                finish booting. In that case, the application code, not RedBoot
                will clear the PCI retry bit."
        }

        cdl_option CYGPKG_HAL_ARM_IQ80310_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the XScale IQ80310 HAL. These flags are used
		in addition to the set of global flags."
        }

        cdl_option CYGPKG_HAL_ARM_IQ80310_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the XScale IQ80310 HAL. These flags are
		removed from the set of global flags if present."
        }

        cdl_option CYGPKG_HAL_ARM_IQ80310_TESTS {
            display "XScale IQ80310 tests"
            flavor  data
            no_define
            calculated { "" }
            description   "
                This option specifies the set of tests for the XScale IQ80310 HAL."
        }
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { CYG_HAL_STARTUP == "RAM" ?       "arm_iq80310_ram" : \
                     CYGSEM_HAL_ARM_IQ80310_ARMBOOT ? "arm_iq80310_roma" : \
	                                              "arm_iq80310_rom" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_iq80310_ram.ldi>" : \
                         CYGSEM_HAL_ARM_IQ80310_ARMBOOT ? "<pkgconf/mlt_arm_iq80310_roma.ldi>" : \
                                                    "<pkgconf/mlt_arm_iq80310_rom.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_iq80310_ram.h>" : \
                         CYGSEM_HAL_ARM_IQ80310_ARMBOOT ? "<pkgconf/mlt_arm_iq80310_roma.h>" : \
                                                    "<pkgconf/mlt_arm_iq80310_rom.h>" }
        }
    }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "ROM" }
        description   "
            Enable this option if this program is to be used as a ROM monitor,
            i.e. applications will be loaded into RAM on the board, and this
            ROM monitor may process exceptions or interrupts generated from the
            application. This enables features such as utilizing a separate
            interrupt stack when exceptions are generated."
    }

    cdl_option CYGSEM_HAL_USE_ROM_MONITOR {
         display       "Work with a ROM monitor"
         flavor        booldata
         legal_values  { "Generic" "GDB_stubs" }
         default_value { CYG_HAL_STARTUP == "RAM" ? "GDB_stubs" : 0 }
         parent        CYGPKG_HAL_ROM_MONITOR
         requires      { CYG_HAL_STARTUP == "RAM" }
         description   "
             Support can be enabled for different varieties of ROM monitor.
             This support changes various eCos semantics such as the encoding
             of diagnostic output, or the overriding of hardware interrupt
             vectors.
             Firstly there is \"Generic\" support which prevents the HAL
             from overriding the hardware vectors that it does not use, to
             instead allow an installed ROM monitor to handle them. This is
             the most basic support which is likely to be common to most
             implementations of ROM monitor.
             \"GDB_stubs\" provides support when GDB stubs are included in
             the ROM monitor or boot ROM."
     }

    cdl_component CYGPKG_REDBOOT_HAL_OPTIONS {
        display       "Redboot HAL options"
        flavor        none
        no_define
        parent        CYGPKG_REDBOOT
        active_if     CYGPKG_REDBOOT
        description   "
            This option lists the target's requirements for a valid Redboot
            configuration."
    
        cdl_option CYGBLD_BUILD_REDBOOT_BIN {
            display       "Build Redboot ROM binary image"
            active_if     CYGBLD_BUILD_REDBOOT
            default_value 1
            no_define
            description "This option enables the conversion of the Redboot ELF
                         image to a binary image suitable for ROM programming."
    
            compile -library=libextras.a diag/diag.c diag/io_utils.c diag/external_timer.c \
				diag/i557_eep.c diag/pci_serv.c diag/interrupts.c          \
				diag/xscale_test.c diag/flash.c diag/cycduart.c            \
                                diag/ether_test.c diag/memtest.c diag/test_menu.c          \
				diag/irq.S
    
            make -priority 325 {
                <PREFIX>/bin/redboot.bin : <PREFIX>/bin/redboot.elf
                $(OBJCOPY) --strip-debug $< $(@:.bin=.img) 
                $(OBJCOPY) -O srec $< $(@:.bin=.srec)
                $(OBJCOPY) -O binary $< $@
            }
        }
    }

}
