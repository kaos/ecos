# ====================================================================
#
#      flash_mbx.cdl
#
#      FLASH memory - Hardware support on Motorola PowerPC/860
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Original data:  gthomas
# Contributors:
# Date:           2000-07-26
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_FLASH_MBX {
    display       "Motorola PowerPC/860 FLASH memory support"

    parent        CYGPKG_IO_FLASH
    active_if	  CYGPKG_IO_FLASH
    requires	  CYGPKG_HAL_POWERPC_MBX

    compile       powerpc_mbx_flash.c

    # Arguably this should do in the generic package
    # but then there is a logic loop so you can never enable it.
    cdl_interface CYGINT_DEVS_FLASH_AMD_AM29XXXXX_REQUIRED {
        display   "Generic AMD AM29F040 driver required"
    }

    implements    CYGINT_DEVS_FLASH_AMD_AM29XXXXX_REQUIRED
    requires      CYGHWR_DEVS_FLASH_AMD_AM29F040B
}
