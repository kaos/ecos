# ====================================================================
#
#      hal_i386_pc.cdl
#
#      PC/i386 target HAL package configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  jskov
# Contributors:
# Date:           1999-11-01
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_I386_PC {
    display  "i386 PC Target"
    parent        CYGPKG_HAL_I386
    define_header hal_i386_pc.h
    include_dir   cyg/hal
    description   "
           The i386 PC Target HAL package provides the 
           support needed to run eCos binaries on an i386 PC."

    compile       hal_diag.c plf_misc.c plf_stub.c

    implements    CYGINT_HAL_DEBUG_GDB_STUBS
    implements    CYGINT_HAL_DEBUG_GDB_STUBS_BREAK
    implements	  CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT
    implements	  CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT_GUARANTEED

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H   <pkgconf/hal_i386.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_i386_pc.h>"
        puts $::cdl_header ""
        puts $::cdl_header "#define HAL_PLATFORM_CPU    \"I386\""
        puts $::cdl_header "#define HAL_PLATFORM_BOARD  \"PC\""
        puts $::cdl_header "#define HAL_PLATFORM_EXTRA  \"\""
	puts $::cdl_header "#include <pkgconf/hal_i386_pcmb.h>"
        puts $::cdl_header ""
    }

    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        legal_values  {"RAM" "FLOPPY" "ROM"}
        default_value {"RAM"}
	no_define
	define -file system.h CYG_HAL_STARTUP
        description   "
            It is possible to configure eCos for the PC target to build for
            RAM startup (generally when being run under an existing
            Monitor program like RedBoot), FLOPPY startup (for writing
            to a floppy disk, which can then be used for booting
            on PCs with a standard BIOS), or ROM startup (for writing
            straight to a boot ROM/Flash). ROM startup is experimental
            at this time."
    }
        
    cdl_option CYGBLD_BUILD_I386_ROMBOOT {
	display       "Build ROM bootstrap code"
	calculated    { CYG_HAL_STARTUP == "ROM" }

	make {
	    <PREFIX>/lib/romboot.ld: <PACKAGE>/src/romboot.ld
	    cp $< $@
	}
	
	make {
	    <PREFIX>/bin/romboot.elf : <PACKAGE>/src/romboot.S
	    @sh -c "mkdir -p $(dir $@)"
	    $(CC) -Wp,-MD,romboot.tmp $(INCLUDE_PATH) -nostdlib -Wl,-static -T$(PREFIX)/lib/romboot.ld -o $@ $<
	    @echo $@ ": \\" > $(notdir $@).deps
	    @tail +2 romboot.tmp >> $(notdir $@).deps
	    @echo >> $(notdir $@).deps
	    @rm romboot.tmp
	}
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD {
        display       "Diagnostic serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 57600 115200
        default_value 38400
        description   "
            This option selects the baud rate used for the diagnostic port.
            Note: this should match the value chosen for the GDB port if the
            diagnostic and GDB port are the same."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_BAUD {
        display       "GDB serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 57600 115200
        default_value 38400
        description   "
            This option controls the baud rate used for the GDB connection."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
        display		"Number of communication channels on the board"
        flavor		data
        legal_values	1 to 3
	default_value	{ CYGSEM_HAL_I386_PC_DIAG_SCREEN ? 3 : 2 }
	description	"
	    This define the number of serial ports that will be used by the HAL.
	    Ports 0 and 1 equate to COM1 and COM2 and port 2 is the PC screen and
	    keyboard."
    }
 
    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
        display          "Debug serial port"
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
            On PCs with two serial ports, this option
            chooses which port will be used to connect to a host
            running GDB."
     }

     cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_DEFAULT {
          display       "Default console channel."
          flavor        data
          legal_values  0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
          default_value 0
     }
 
     cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
         display          "Diagnostic serial port"
         flavor data
         legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
         default_value    CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_DEFAULT
         description      "
            On PCs with two serial ports, this option
            chooses which port will be used for diagnostic output.
	    Selecting port 2 will cause the PC screen to be used."
     }

     cdl_option CYGSEM_HAL_I386_PC_DIAG_SCREEN {
	 display       "Output to PC screen"
	 flavor        bool
	 default_value 1
	 implements CYGINT_HAL_I386_PCMB_SCREEN_SUPPORT
	 description "This option enables use of the PC screen and keyboard as a
	             third virtual serial device."
     }
     
    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        parent  CYGPKG_NONE
        description   "
	    Global build options including control over
	    compiler flags, linker flags and choice of toolchain."


        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "i386-elf" }
            description "
                This option specifies the command prefix used when
                invoking the build tools. If your host operating system
                is Linux you can set this to empty to use your native tools.
                If so, your native gcc must be gcc-2.95.2 or later, and
                \"ld -v\" must report a version more recent than 2.9.1."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { "-Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority" }
            description   "
                This option controls the global compiler flags which
                are used to compile all packages by
                default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { "-g -nostdlib -Wl,--gc-sections -Wl,-static" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }

        cdl_option CYGBLD_BUILD_GDB_STUBS {
            display "Build GDB stub loader image"
            default_value 0
            requires { CYG_HAL_STARTUP == "FLOPPY" }
            requires CYGSEM_HAL_ROM_MONITOR
            requires CYGBLD_BUILD_COMMON_GDB_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
            requires ! CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT
            requires ! CYGDBG_HAL_DEBUG_GDB_CTRLC_SUPPORT
            requires ! CYGDBG_HAL_DEBUG_GDB_THREAD_SUPPORT
            requires ! CYGDBG_HAL_COMMON_INTERRUPTS_SAVE_MINIMUM_CONTEXT
            requires ! CYGDBG_HAL_COMMON_CONTEXT_SAVE_MINIMUM
            no_define
            description "
                This option enables the building of the GDB stubs for the
                board. The common HAL controls takes care of most of the
                build process, but the final conversion from ELF image to
                binary data is handled by the platform CDL, allowing
                relocation of the data if necessary."

            make -priority 320 {
                <PREFIX>/bin/gdb_module.bin : <PREFIX>/bin/gdb_module.img
                $(OBJCOPY) -O binary $< $@
            }
        }
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { CYG_HAL_STARTUP == "RAM" ? "i386_pc_ram" : \
		     CYG_HAL_STARTUP == "ROM" ? "i386_pc_rom" : \
	                                        "i386_pc_floppy" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_i386_pc_ram.ldi>" : \
		         CYG_HAL_STARTUP == "ROM" ? "<pkgconf/mlt_i386_pc_rom.ldi>" : \
                                                    "<pkgconf/mlt_i386_pc_floppy.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_i386_pc_ram.h>" : \
		         CYG_HAL_STARTUP == "ROM" ? "<pkgconf/mlt_i386_pc_rom.h>" : \
                                                    "<pkgconf/mlt_i386_pc_floppy.h>" }
        }
    }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
	
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "FLOPPY" || CYG_HAL_STARTUP == "ROM" }
	requires      { !CYGHWR_HAL_I386_FPU_SWITCH_LAZY }
        description   "
            Enable this option if this program is to be used as a ROM monitor,
            i.e. applications will be loaded into RAM on the board, and this
            ROM monitor may process exceptions or interrupts generated from the
            application. This enables features such as utilizing a separate
            interrupt stack when exceptions are generated."
    }

    cdl_option CYGSEM_HAL_USE_ROM_MONITOR {
         display       "Work with a ROM monitor"
         flavor        booldata
         legal_values  { "Generic" "GDB_stubs" }
         default_value { CYG_HAL_STARTUP == "RAM" ? "GDB_stubs" : 0 }
         parent        CYGPKG_HAL_ROM_MONITOR
         requires      { CYG_HAL_STARTUP == "RAM" }
         description   "
             Support can be enabled for different varieties of ROM monitor.
             This support changes various eCos semantics such as the encoding
             of diagnostic output, or the overriding of hardware interrupt
             vectors.
             Firstly there is \"Generic\" support which prevents the HAL
             from overriding the hardware vectors that it does not use, to
             instead allow an installed ROM monitor to handle them. This is
             the most basic support which is likely to be common to most
             implementations of ROM monitor.
             \"GDB_stubs\" provides support when GDB stubs are included in
             the ROM monitor or boot ROM."
     }

    cdl_component CYGPKG_REDBOOT_HAL_OPTIONS {
        display       "Redboot HAL options"
        flavor        none
        no_define
        parent        CYGPKG_REDBOOT
        active_if     CYGPKG_REDBOOT
        description   "
            This option lists the target's requirements for a valid Redboot
            configuration."
    
        cdl_component CYGBLD_BUILD_REDBOOT_BIN {
            display       "Build RedBoot binary image"
            no_define
            default_value 1

            cdl_option CYGBLD_BUILD_REDBOOT_BIN_FLOPPY {
                display       "Build Redboot FLOPPY binary image"
                active_if     CYGBLD_BUILD_REDBOOT
                active_if     { CYG_HAL_STARTUP == "FLOPPY" }
                calculated    1
                no_define
                description "This option enables the conversion of the Redboot 
                             ELF image to a binary image suitable for
                             copying to a floppy disk."
        
                make -priority 325 {
                    <PREFIX>/bin/redboot.bin : <PREFIX>/bin/redboot.elf
                    $(OBJCOPY) -O binary $< $@
                }
            }
    
            cdl_option CYGBLD_BUILD_REDBOOT_BIN_ROM {
                display       "Build Redboot ROM binary image"
                active_if     CYGBLD_BUILD_REDBOOT
                active_if     { CYG_HAL_STARTUP == "ROM" }
                calculated    1
                no_define
                description "This option enables the conversion of the Redboot
                             ELF image to a binary image suitable for ROM
                             programming."
                
                make -priority 325 {
                    <PREFIX>/bin/redboot.bin : <PREFIX>/bin/redboot.elf
                    $(OBJCOPY) -O binary $< $(@:.bin=.img)
                    $(OBJCOPY) -O binary $(PREFIX)/bin/romboot.elf $(PREFIX)/bin/romboot.img
                    dd if=/dev/zero of=$@ bs=1024 count=64 conv=sync
                    dd if=$(@:.bin=.img) of=$@ bs=512 conv=notrunc,sync
                    dd if=$(PREFIX)/bin/romboot.img of=$@ bs=256 count=1 seek=255 conv=notrunc
                }
            }
        }            
    }     
}

