# ====================================================================
#
#      compat.cdl
#
#      Maths library compatibility related configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  jlarmour
# Contributors:
# Date:           1999-07-07
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_interface CYGINT_LIBM_COMPAT {
    requires 1 == CYGINT_LIBM_COMPAT
}

cdl_option CYGSEM_LIBM_COMPAT_IEEE_ONLY {
    display       "IEEE-only"
    default_value 0
    implements    CYGINT_LIBM_COMPAT
    description   "
        The math library can be hard-coded to only
        behave in one compatibility mode - IEEE. This
        cannot be changed at run-time. IEEE mode is the
        most minimal of the compatibility modes, and so
        this will best help code size and speed, as well
        as omitting the code for other compatibility
        modes. If not defined, the math library can be
        set at run-time to any of the supported
        compatibility modes."
}

cdl_component CYGNUM_LIBM_COMPATIBILITY {
    display       "Default mode"
    flavor        booldata
    requires      CYGPKG_LIBC
    implements    CYGINT_LIBM_COMPAT
    legal_values  { "POSIX" "IEEE" "XOPEN" "SVID" }
    default_value { "POSIX" }
    define        CYGPKG_LIBM_COMPATIBILITY_DEFAULT
    description   "
        If you want to have support for more than one
        compatibility mode settable at run-time, rather
        than hard-coded IEEE mode, this component lets
        you choose which mode should be the default."

    cdl_option CYGNUM_LIBM_COMPAT_DEFAULT {
      	display       "Numeric representation"
	flavor        data
	calculated   { \
            CYGNUM_LIBM_COMPATIBILITY == "POSIX" ? "CYGNUM_LIBM_COMPAT_POSIX" :\
            CYGNUM_LIBM_COMPATIBILITY == "IEEE"  ? "CYGNUM_LIBM_COMPAT_IEEE" :\
            CYGNUM_LIBM_COMPATIBILITY == "XOPEN" ? "CYGNUM_LIBM_COMPAT_XOPEN" :\
            CYGNUM_LIBM_COMPATIBILITY == "SVID"  ? "CYGNUM_LIBM_COMPAT_SVID" :\
	    "<undefined>" \
        }
	description	"
	    This option automatically defines the default compatibility
	    mode for numeric representation in terms of the values used
	    to set that mode at run-time."
    }
}

cdl_option CYGFUN_LIBM_SVID3_scalb {
    display       "SVID3-style scalb()"
    default_value 1
    description   "
        SVID3 defined the scalb() function as double
        scalb(double, double) rather than double
        scalb(double, int) which is used by IBM, DEC, and
        probably others. Enabling this option chooses
        the (double, double) version. Note there is a
        function double scalbn(double, int) which is
        unaffected by this choice."
}

cdl_option CYGSYM_LIBM_NO_XOPEN_SVID_NAMESPACE_POLLUTION {
    display       "Reduce namespace pollution"
    default_value 0
    description   "
        If you do not want to use either the X/Open or
        SVID3 compatibility modes, you may want to define
        this option to reduce the chance of namespace
        pollution. This is particularly likely to occur
        here as these standards define symbols with
        names that often appear in applications, such as
        exception, DOMAIN, OVERFLOW, etc. If your
        application also used these names, it may cause
        problems."
}

cdl_option CYGSEM_LIBM_USE_STDERR {
    display       "Output to stderr for math errors"
    requires      !CYGSEM_LIBM_COMPAT_IEEE_ONLY
    requires      CYGPKG_LIBC_STDIO
    default_value 0
    description   "
        The SVID3 standard says that error
        messages should be output on the stderr console
        output stream. This option allows this ability
        to be explicitly controlled. However, this still
        only has an effect in SVID3 compatibility mode."
}
