# ====================================================================
#
#      usbs_eth.cdl
#
#      USB slave-side ethernet package.
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000, 2001 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      bartv
# Original data:  bartv
# Contributors:
# Date:           2000-10-04
#
#####DESCRIPTIONEND####
# ====================================================================

cdl_package CYGPKG_IO_USB_SLAVE_ETH {
    display     "USB slave ethernet support"
    include_dir "cyg/io/usb"
    parent      CYGPKG_IO_USB_SLAVE
    requires    { CYGHWR_IO_USB_SLAVE_OUT_ENDPOINTS >= 1 }
    requires    { CYGHWR_IO_USB_SLAVE_IN_ENDPOINTS >= 1 }
    compile     usbseth.c
    implements  CYGINT_IO_USB_SLAVE_CLIENTS
    doc         io-usb-slave-eth.html
    
    description "
        The USB slave ethernet package supports the development
        of USB peripherals which provide an ethernet service to
        the host machine. Such a peripheral could be a simple
        USB-ethernet converter, or it could be rather more
        complicated internally."

    cdl_component CYGPKG_USBS_ETHDRV {
	display         "Provide a driver for a TCP/IP stack."
        requires        CYGPKG_IO_ETH_DRIVERS
	implements      CYGHWR_NET_DRIVERS
	default_value   CYGPKG_NET
	compile         -library=libextras.a usbsethdrv.c

	description "
	    The primary purpose of USB slave ethernet support is to provide
	    an ethernet service to the USB host. This is very different
	    from a conventional network driver which provides a service
            to a TCP/IP stack running inside the peripheral. If this
	    component is enabled then the USB-ethernet code will implement
	    an eCos network driver, thus supporting both a host-side TCP/IP
	    stack and an eCos stack. This raises issues such as enabling
	    the bridge code in the stack, and the package documentation
            should be consulted for further information."

	cdl_option CYGFUN_USBS_ETHDRV_STATISTICS {
	    display       "Maintain traffic statistics"
	    flavor        bool
	    default_value CYGPKG_SNMPAGENT
	    description "
	        The USB network device driver can maintain some statistics
                about traffic, for example the number of incoming and
	        outgoing packets. These statistics are intended mainly
	        for SNMP agent software."
	}

	cdl_option CYGDAT_USBS_ETHDRV_NAME {
	    display       "Name to use for this network device"
	    flavor        data
	    default_value { "\"eth0\"" }
	    description "
	        The name of this network device for control purposes.
	    "
	}

	cdl_option CYGPRI_USBS_ETHDRV_ETH0 {
	    display       "Enable/disable generic eth0 configury"
	    flavor        bool
	    calculated    { "\"eth0\"" == CYGDAT_USBS_ETHDRV_NAME }
	    implements    CYGHWR_NET_DRIVER_ETH0
	}
	cdl_option CYGPRI_USBS_ETHDRV_ETH1 {
	    display       "Enable/disable generic eth1 configury"
	    flavor        bool
	    calculated    { "\"eth1\"" == CYGDAT_USBS_ETHDRV_NAME }
	    implements    CYGHWR_NET_DRIVER_ETH1
	}
    }
}
