# ====================================================================
#
#      semas.cdl
#
#      uITRON semaphore related configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  hmt
# Contributors:
# Date:           1999-07-07
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_option CYGNUM_UITRON_SEMAS {
    display       "Number of semaphores"
    flavor        data
    legal_values  1 to 65535
    default_value 3
    description   "
        The number of uITRON semaphores present in the system.
        Valid semaphore object IDs will range from 1 to this value."
}
cdl_component CYGPKG_UITRON_SEMAS_CREATE_DELETE {
    display       "Support create and delete"
    flavor        bool
    default_value 1
    description   "
        Support semaphore create and delete operations (cre_sem, del_sem).
        Otherwise all semaphores are created, up to the number specified 
        above."

    cdl_option CYGNUM_UITRON_SEMAS_INITIALLY {
        display       "Number of semaphores created initially"
        flavor        data
        legal_values  0 to 65535
        default_value 3
        description   "
            The number of uITRON semaphores initially created.
            This number should not be more than the number
            of semaphores in the system, though setting it to a large
            value to mean 'all' is acceptable.
            Initially, only semaphores numbered 1 to this number exist;
            higher numbered ones must be created before use.
            It is only useful to initialize semaphores up to this number;
            higher numbered ones must be created in order to use them,
            and so they will be re-initialized."
    }
}
cdl_component CYGPKG_UITRON_SEMAS_ARE_INITIALIZED {
    display       "Initialize semaphore counts"
    flavor        bool
    default_value 0
    description   "
        Initialize semaphores to specific count values.
        Otherwise semaphores are initialized with the count
        set to zero."

    cdl_option CYGDAT_UITRON_SEMA_INITIALIZERS {
        display       "Static initializers"
        parent        CYGPKG_UITRON_SEMAS_ARE_INITIALIZED
        flavor        data
        default_value {"CYG_UIT_SEMA(  0 ),\
                        CYG_UIT_SEMA(  0 ),\
                        CYG_UIT_SEMA(  0 )"}
        description   "
            A list of initializers separated by commas,
            one per line.
            An initializer is 'CYG_UIT_SEMA(INITIAL-COUNT)'
            or 'CYG_UIT_SEMA_NOEXS' for slots above the number
            initially to be created, when create and delete
            operations are supported.
            Note: this option is invoked in the context of a
            C++ array initializer, between curly brackets.
            Ensure that the number of initializers here exactly
            matches the total number of semaphores specified."
    }
}
