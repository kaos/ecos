# ====================================================================
#
#      v85x_edb_v850_disk.cdl
#
#      Elatec v850 development board disk package.
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 2003 Savin Zlobec 
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      savin
# Contributors:
# Date:           2003-08-21
#
#####DESCRIPTIONEND####
# ====================================================================

cdl_package CYGPKG_DEVS_DISK_V85X_EDB_V850 {
    display     "Disk driver for Elatec v850 development board"
    
    parent      CYGPKG_IO_DISK_DEVICES
    active_if   CYGPKG_IO_DISK
    active_if   CYGPKG_HAL_V85X_EDB_V850

    compile     -library=libextras.a   v85x_edb_v850_disk.c
    
    cdl_component CYGVAR_DEVS_DISK_V85X_EDB_V850_DISK0 {
    	display         "Provide disk 0 device"
        flavor          bool
        default_value   0
        description     "Elatec v850 development board disk 0 driver."
        
        cdl_option CYGDAT_IO_DISK_V85X_EDB_V850_DISK0_NAME {
            display       "Device name for disk 0 device"
            flavor        data
            default_value {"\"/dev/v85xdisk0/\""}
        }
    }
}

# EOF v85x_edb_v850_disk.cdl
