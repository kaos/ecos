# ====================================================================
#
#      hal_powerpc.cdl
#
#      PowerPC architectural HAL package configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  bartv
# Contributors:
# Date:           1999-11-02
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_POWERPC {
    display  "PowerPC architecture"
    parent        CYGPKG_HAL
    hardware
    include_dir   cyg/hal
    define_header hal_powerpc.h
    description   "
        The PowerPC architecture HAL package provides generic
        support for this processor architecture. It is also
        necessary to select a specific target platform HAL
        package."

    cdl_interface CYGINT_HAL_POWERPC_VARIANT {
        display  "Number of variant implementations in this configuration"
        no_define
        requires 1 == CYGINT_HAL_POWERPC_VARIANT
    }

    compile       hal_misc.c context.S ppc_stub.c hal_intr.c

    # The "-o file" is a workaround for CR100958 - without it the
    # output file would end up in the source directory under CygWin.
    # n.b. grep does not behave itself under win32
    make -priority 1 {
        <PREFIX>/include/cyg/hal/ppc_offsets.inc : <PACKAGE>/src/hal_mk_defs.c
        $(CC) $(CFLAGS) $(INCLUDE_PATH) -Wp,-MD,ppc_offsets.tmp -o hal_mk_defs.tmp -S $<
        fgrep .equ hal_mk_defs.tmp | sed s/#// > $@
        @echo $@ ": \\" > $(notdir $@).deps
        @tail -n +2 ppc_offsets.tmp >> $(notdir $@).deps
        @echo >> $(notdir $@).deps
        @rm ppc_offsets.tmp hal_mk_defs.tmp
    }

    make {
        <PREFIX>/lib/vectors.o : <PACKAGE>/src/vectors.S
        $(CC) -Wp,-MD,vectors.tmp $(INCLUDE_PATH) $(CFLAGS) -c -o $@ $<
        @echo $@ ": \\" > $(notdir $@).deps
        @tail -n +2 vectors.tmp >> $(notdir $@).deps
        @echo >> $(notdir $@).deps
        @rm vectors.tmp
    }

    make {
        <PREFIX>/lib/target.ld: <PACKAGE>/src/powerpc.ld
        $(CC) -E -P -Wp,-MD,target.tmp -DEXTRAS=1 -xc $(INCLUDE_PATH) $(CFLAGS) -o $@ $<
        @echo $@ ": \\" > $(notdir $@).deps
        @tail -n +2 target.tmp >> $(notdir $@).deps
        @echo >> $(notdir $@).deps
        @rm target.tmp
    }

    cdl_option CYGSEM_HAL_POWERPC_RESET_USES_JUMP {
        display       "RESET vector jumps to startup"
        default_value 0
        description   "
            Some platforms may need this for ROMRAM startup."
    }

    cdl_option CYGSEM_HAL_POWERPC_COPY_VECTORS {
        display       "Copy exception vectors to RAM"
        default_value { (CYG_HAL_STARTUP != "RAM" ||
                         CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS) ? 1 : 0 }
        requires      ! CYGSEM_HAL_USE_ROM_MONITOR
        description   "
            Enable this option to force exception vectors to be copied
            to the vector base on startup. For RAM startup this is normally
            disabled since the vectors would already have been provided
            by the GDB stubs - but it's possible to override, thus taking
            full control of the target. For ROM startup it is desirable to
            enable this option if the vector base is set to RAM since
            accessing vectors in ROM is normally slower. But if memory is
            tight the vectors can be left in ROM."
    }

    cdl_option CYGHWR_HAL_POWERPC_NEED_VECTORS {
        display       "Exception vectors inclusion"
        description   "
            If eCos can rely on the target environment to provide
            eCos compatible vector code, there is no reason to include
            the additional data in application images. This option controls
            the inclusion of the vector code."
        # Platform HALs and startup configuration controls this setting.
        calculated { ((CYGHWR_HAL_POWERPC_FORCE_VECTORS ||
                       CYG_HAL_STARTUP != "RAM" ||
                       CYGSEM_HAL_POWERPC_COPY_VECTORS) &&
                      ! CYGSEM_HAL_USE_ROM_MONITOR)
                      ? 1 : 0 }
    }

    cdl_option CYGHWR_HAL_POWERPC_VECTOR_BASE {
        display       "Exception vectors location"
        description   "
            PowerPC exception vectors can reside either at 0x00000000 or
            0xfff00000. The startup type and platform HAL controls which
            is used."
        flavor        data
        calculated { (! CYGHWR_HAL_POWERPC_FORCE_VECTOR_BASE_LOW && 
                       (CYGHWR_HAL_POWERPC_FORCE_VECTOR_BASE_HIGH ||
                       (CYG_HAL_STARTUP != "RAM" &&
                        ! CYGSEM_HAL_POWERPC_COPY_VECTORS)))
                      ? 0xfff00000 : 0x00000000 }
    }

    cdl_option CYGHWR_HAL_POWERPC_ENABLE_MMU {
        display       "Enable MMU"
        default_value { !CYGHWR_HAL_POWERPC_DISABLE_MMU }
        description   "
            Some platforms do not want the MMU enabled."
    }

    cdl_option CYGDBG_HAL_POWERPC_FRAME_WALLS {
        display       "Exception stack-frame walls"
        default_value 0
        description   "
            Enable this option to put \"walls\" around the exception
            frames. This can ease analyzing the stack contents when
            debugging."
    }

    cdl_option CYGSEM_REDBOOT_HAL_LINUX_BOOT {
        active_if      { CYGSEM_REDBOOT_PLF_LINUX_BOOT == 1 }
        display        "Support booting Linux via RedBoot"
        flavor         bool
        default_value  1
        description    "
           This option enables RedBoot to support booting of a Linux kernel."

        compile -library=libextras.a redboot_linux_exec.c
    }

    cdl_component CYGPKG_HAL_POWERPC_OPTIONS {
        display "PowerPC build options"
        flavor  none
        no_define
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_HAL_POWERPC_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the PowerPC HAL. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_HAL_POWERPC_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the PowerPC HAL. These flags are removed from
                the set of global flags if present."
        }

        cdl_option CYGPKG_HAL_POWERPC_TESTS {
            display "PowerPC tests"
            flavor  data
            no_define
            calculated { "" }
            description   "
                This option specifies the set of tests for the PowerPC HAL."
        }
    }

    cdl_option CYGBLD_LINKER_SCRIPT {
        display "Linker script"
        flavor data
	no_define
        calculated  { "src/powerpc.ld" }
    }
}
