# ====================================================================
#
#	davicom_dm9000_eth_drivers.cdl
#
#	Davicom dm9000 ethernet driver
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2003, 2004 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      msalter
# Original data:
# Contributors:
# Date:           2004-3-18
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_DAVICOM_DM9000 {
    display       "Davicom DM9000 ethernet driver"
    description   "Ethernet driver for Davicom DM9000 NIC."

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if     CYGPKG_IO_ETH_DRIVERS

    active_if     CYGINT_DEVS_ETH_DAVICOM_DM9000_REQUIRED

    define_proc {
        puts $::cdl_header "#include CYGDAT_DEVS_ETH_DAVICOM_DM9000_CFG";
    }

    compile       -library=libextras.a if_dm9000.c

    cdl_option CYGSEM_DEVS_ETH_DAVICOM_DM9000_WRITE_EEPROM {
        display "SIOCSIFHWADDR records ESA (MAC address) in EEPROM"
        default_value 0
        description   "
            The ioctl() socket call with operand SIOCSIFHWADDR sets the
            interface hardware address - the MAC address or Ethernet Station
            Address (ESA).  This option causes the new MAC address to be
            written into the EEPROM associated with the interface, so that the
            new MAC address is permanently recorded.  Doing this should be a
            carefully chosen decision, hence this option."
    }

    cdl_option CYGNUM_DEVS_ETH_DAVICOM_DM9000_DEV_COUNT {
	display "Number of supported interfaces."
	calculated    { CYGINT_DEVS_ETH_DAVICOM_DM9000_REQUIRED }
        flavor        data
	description   "
	    This option selects the number of PCMCIA cards to
            be supported by the driver."
    }

    cdl_component CYGPKG_DEVS_ETH_DAVICOM_DM9000_OPTIONS {
        display "Davicom dm9000 ethernet driver build options"
        flavor  none
	no_define

        cdl_option CYGPKG_DEVS_ETH_DAVICOM_DM9000_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the Davicom DM9000 ethernet driver package.
                These flags are used in addition to the set of
                global flags."
        }
    }
}
# EOF davicom_dm9000_eth_drivers.cdl
