# ====================================================================
#
#      hal_h8300_h8s.cdl
#
#      H8S variant architectural HAL package configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      ysato
# Original data:  nickg
# Contributors:   ysato
# Date:           2003-01-01
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_H8300_H8S {
    display "H8S variant"
    parent        CYGPKG_HAL_H8300
    implements CYGINT_HAL_H8300_VARIANT
    hardware
    include_dir   cyg/hal
    define_header hal_h8300_h8s.h
    description   "
           The H8S variant HAL package provides generic
           support for this processor architecture. It is also
           necessary to select a specific target platform HAL
           package."

    define_proc {
        puts $::cdl_header "#include <pkgconf/hal_h8300.h>"
    }

    compile       var_misc.c h8s_stub.c

    make {
        <PREFIX>/lib/target.ld: <PACKAGE>/src/h8300_h8s.ld
        $(CC) -E -P -Wp,-MD,target.tmp -DEXTRAS=1 -xc $(INCLUDE_PATH) $(CFLAGS) -o $@ $<
        @echo $@ ": \\" > $(notdir $@).deps
        @tail +2 target.tmp >> $(notdir $@).deps
        @echo >> $(notdir $@).deps
        @rm target.tmp
    }

    cdl_option CYGBLD_LINKER_SCRIPT {
        display "Linker script"
        flavor data
	no_define
        calculated  { "src/h8300_h8s.ld" }
    }

    cdl_component CYGHWR_HAL_H8S_CLOCK_SETTINGS {
        display          "H8S on-chip generic clock controls"
        description      "
            The various clocks used by the system are controlled by
            these options, some of which are derived from platform
            settings."
        flavor        none
        no_define

 	cdl_option CYGHWR_HAL_H8300_DIVIDER_RATE {
 	    display	     "Divider Rate (1/n)"
 	    flavor	     data
             legal_values     { 1 2 4 8 }
 	    default_value    1
 	    description	     "
               The system clock divide rate setting"
 	}
 	cdl_option CYGHWR_HAL_H8300_MULT_RATE {
 	    display	     "PLL Multiplier Rate (Nx)"
 	    flavor	     data
             legal_values     { 1 2 4 }
 	    default_value    1
 	    description	     "
               The system clock divide rate setting"
 	}
        cdl_option CYGHWR_HAL_H8300_PROCESSOR_SPEED {
             display          "Processor clock speed (MHz)"
             flavor           data
             calculated       { CYGHWR_HAL_H8300_CPG_INPUT * CYGHWR_HAL_H8300_MULT_RATE / CYGHWR_HAL_H8300_DIVIDER_RATE }
             description      "
                 The core (CPU) speed is computed from
                 the input clock speed and the divider setting."
         }
    }
}
