# ====================================================================
#
#      synch.cdl
#
#      configuration data related to the kernel synchronization primitives
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  nickg
# Contributors:
# Date:           1999-07-05
#
#####DESCRIPTIONEND####
#
# ====================================================================


cdl_component CYGSEM_KERNEL_SYNCH_MUTEX_PRIORITY_INVERSION_PROTOCOL {
    display      "Priority inversion protection protocols"
    flavor       booldata
    legal_values { "SIMPLE" }
    default_value { "SIMPLE" }
    active_if    { CYGSEM_KERNEL_SCHED_MLQUEUE }
    requires     { CYGINT_KERNEL_SCHEDULER_UNIQUE_PRIORITIES == 0 }
    description "
        This component controls the protocols used to protect mutexes against
        priority inversion. If this option is enabled it defines which
        algorithm is used to implement this protection. At present only
        one such algorithm is defined: \"SIMPLE\". The implementation
        will only work in the mlqueue scheduler, and it does not handle the
        rare case of nested mutexes completely correctly. However it is
        both fast and deterministic."

    cdl_option  CYGSEM_KERNEL_SYNCH_MUTEX_PRIORITY_INVERSION_PROTOCOL_INHERIT {
	display       "Enable priority inheritance protocol"
	default_value 1
	implements CYGINT_KERNEL_SYNCH_MUTEX_PRIORITY_INVERSION_PROTOCOL_COUNT
	description   "
	    This option enables priority inheritance protocol. This protocol
	    causes the owner of a mutex to be executed at the highest priority
	    of the threads waiting for access to the mutex."
    }

    cdl_option CYGSEM_KERNEL_SYNCH_MUTEX_PRIORITY_INVERSION_PROTOCOL_CEILING {
	display       "Enable priority ceiling protocol"
	default_value 1
	implements CYGINT_KERNEL_SYNCH_MUTEX_PRIORITY_INVERSION_PROTOCOL_COUNT	
	description   "
	    This option enables priority ceiling protocol. This protocol
	    causes the owner of a mutex to be executed at a  priority
	    associated with the mutex."
    }

    cdl_option CYGSEM_KERNEL_SYNCH_MUTEX_PRIORITY_INVERSION_PROTOCOL_NONE {
	display       "No priority inversion protocol"
	default_value 1
	implements CYGINT_KERNEL_SYNCH_MUTEX_PRIORITY_INVERSION_PROTOCOL_COUNT	
	description   "
	    This option enables the ability to have no priority inversion protocol.
	    It is equivalent to disabling the priority inversion protocol at
	    the top level, but is necessary for the runtime and default
	    selection options."
    }

    cdl_option CYGSEM_KERNEL_SYNCH_MUTEX_PRIORITY_INVERSION_PROTOCOL_DEFAULT {
	display      "Default priority inversion protocol"
	flavor       data
	legal_values { "INHERIT" "CEILING" "NONE" }
	default_value { CYGSEM_KERNEL_SYNCH_MUTEX_PRIORITY_INVERSION_PROTOCOL_INHERIT ?
                        "INHERIT" :
                        CYGSEM_KERNEL_SYNCH_MUTEX_PRIORITY_INVERSION_PROTOCOL_CEILING ?
                        "CEILING" : "NONE" }
	description   "
	    This option defines the default inversion protocol used for mutexes that
	    are created without an explicit protocol being specified. The protocol
	    chosen by default is to use priority inheritance if it is present otherwise
	    priority ceiling, or none if neither is present."
    }

    cdl_option CYGSEM_KERNEL_SYNCH_MUTEX_PRIORITY_INVERSION_PROTOCOL_DEFAULT_PRIORITY {
	display       "Default priority ceiling"
	flavor        data
	legal_values  0 to { CYGNUM_KERNEL_SCHED_PRIORITIES - 1 }
	default_value 0
	active_if     { CYGSEM_KERNEL_SYNCH_MUTEX_PRIORITY_INVERSION_PROTOCOL_DEFAULT == "CEILING" }
	description   "
	    This option defines the default priority ceiling to be
	    used if the chosen default priority inversion protocol is
	    priority ceiling protocol. The default value for this is zero,
	    making all such mutexes boost threads to the maximum priority."
    }

    cdl_option CYGSEM_KERNEL_SYNCH_MUTEX_PRIORITY_INVERSION_PROTOCOL_DYNAMIC {
	display        "Specify mutex priority inversion protocol at runtime"
	default_value  1
	active_if      { CYGINT_KERNEL_SYNCH_MUTEX_PRIORITY_INVERSION_PROTOCOL_COUNT > 1 }
	description    "
	    This option controls whether the priority inversion protocol used by
	    a mutex can be specified when that mutex is created."
    }
    
    cdl_interface CYGINT_KERNEL_SYNCH_MUTEX_PRIORITY_INVERSION_PROTOCOL_COUNT {
	display      "Number of protocols selected"
    }
    
}

cdl_option CYGMFN_KERNEL_SYNCH_MBOXT_PUT_CAN_WAIT {
    display       "Message box blocking put support"
    default_value 1
    description   "
        Message boxes can support three different versions of the
        put-message operation. The first is tryput(), which will fail
        if the message box is already full. The other two are the
        ordinary put() function which will block if the message box
        is full, and a timed put() operation which will block for
        upto a certain length of time if the message box is currently
        full. The blocking versions require extra memory in the
        message box data structure and extra code in the other
        message box functions, so they can be disabled if the
        application does not require them. If this option is enabled
        then the system will always provide the blocking put()
        function, and it will also provide the timed put() function
        if thread timers are enabled."
}

cdl_option CYGNUM_KERNEL_SYNCH_MBOX_QUEUE_SIZE {
    display       "Message box queue size"
    flavor        data
    legal_values  1 to 65535
    default_value 10
    description   "
        This configuration option controls the number of messages
        that can be queued in a message box before a non-blocking
        put() operation will fail or a blocking put() operation will
        block. The cost in memory is one pointer per message box for
        each possible message."
}

cdl_option CYGMFN_KERNEL_SYNCH_CONDVAR_TIMED_WAIT {
    display       "Condition variable timed-wait support"
    requires      CYGFUN_KERNEL_THREADS_TIMER
    default_value 1
    description   "
        This option enables the condition variable timed wait
        facility."
}

cdl_option CYGMFN_KERNEL_SYNCH_CONDVAR_WAIT_MUTEX {
    display       "Condition variable explicit mutex wait support"
    default_value 1
    description   "
        This option enables the condition variable explicit mutex wait
        facility. By default condition variables in eCos are created with
        a statically associated mutex. This option permits wait (and timed wait
        if CYGMFN_KERNEL_SYNCH_CONDVAR_TIMED_WAIT is enabled) to provide a
        different mutex as an argument. This makes no difference to the semantics
        the wait operation except that a different mutex will be used during it."
}
