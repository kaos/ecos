# ====================================================================
#
#      hal_arm_sa11x0.cdl
#
#      ARM SA11x0 architectural HAL package configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000, 2001 Red Hat, Inc.
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Original data:  gthomas
# Contributors:
# Date:           2000-05-08
#
#####DESCRIPTIONEND####
#
# ====================================================================
cdl_package CYGPKG_HAL_ARM_SA11X0 {
    display       "ARM SA11X0 architecture"
    parent        CYGPKG_HAL_ARM
    hardware
    include_dir   cyg/hal
    define_header hal_arm_sa11x0.h
    description   "
        This HAL variant package provides generic
        support for the Intel StrongARM SA11x0 processors. It is also
        necessary to select a specific target platform HAL
        package."

    # Let the architectural HAL see this variant's interrupts file -
    # the SA11x0 has no variation between targets here.
    define_proc {
        puts $::cdl_header \
       "#define CYGBLD_HAL_VAR_INTS_H <cyg/hal/hal_var_ints.h>"
    }

    compile       hal_diag.c sa11x0_misc.c

    cdl_option CYGHWR_HAL_ARM_SA11X0_PROCESSOR_CLOCK {
        display       "Processor clock rate"
        active_if     { CYG_HAL_STARTUP == "ROM" }
        flavor        data
        legal_values  59000 73700 88500 103200 118000 132700 147500 162200 176900 191700 206400 221200
        default_value { CYGHWR_HAL_ARM_SA11X0_PROCESSOR_CLOCK_OVERRIDE_DEFAULT ?
                        CYGHWR_HAL_ARM_SA11X0_PROCESSOR_CLOCK_OVERRIDE_DEFAULT : 221200}
        description   "
           The SA-1100 processor can run at various frequencies.
           These values are expressed in KHz.  Note that there are
           several steppings of the SA-1100 rated to run at different
           maximum frequencies.  Check the specs to make sure that your
           particular processor can run at the rate you select here."
    }

    # Real-time clock/counter specifics
    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants"
        flavor        none
        no_define
    
        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            calculated    1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            default_value 100
            description   "
              This option selects the heartbeat rate for the real-time clock.
              The rate is specified in ticks per second.  Change this value
              with caution - too high and your system will become saturated
              just handling clock interrupts, too low and some operations
              such as thread scheduling may become sluggish."
        }
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
            calculated    (3686400/CYGNUM_HAL_RTC_DENOMINATOR)        ;# Clock for OS Timer is 3.6864MHz
        }
    }

    # Control over hardware layout.  
    cdl_interface     CYGHWR_HAL_ARM_SA11X0_UART1 {
        display   "UART1 available as diagnostic/debug channel"
        description "
	  The SA11x0 chip has multiple serial channels which may be
          used for different things on different platforms.  This
          interface allows a platform to indicate that the specified
          serial port can be used as a diagnostic and/or debug channel."
    }

    cdl_interface     CYGHWR_HAL_ARM_SA11X0_UART3 {
        display   "UART3 available as diagnostic/debug channel"
        description "
	  The SA11x0 chip has multiple serial channels which may be
          used for different things on different platforms.  This
          interface allows a platform to indicate that the specified
          serial port can be used as a diagnostic and/or debug channel."
    }

    cdl_option CYGPKG_HAL_ARM_SA11X0_TESTS {
	display "SA11x0 HAL tests"
	flavor  data
	no_define
	calculated { "tests/mmap_test" }
	description   "
	This option specifies the set of tests for the SA11x0 HAL."
    }

    cdl_component CYGPKG_REDBOOT_SA11X0_OPTIONS {
        display       "Redboot for SA11x0 options"
        flavor        none
        no_define
        parent        CYGPKG_REDBOOT
        active_if     CYGPKG_REDBOOT
        description   "
            This option lists the target's requirements for a valid Redboot
            configuration."

        cdl_option CYGSEM_REDBOOT_SA11X0_LINUX_BOOT {
            display        "Support booting Linux via RedBoot"
            flavor         bool
            default_value  1
            description    "
               This option enables RedBoot to support booting of a Linux kernel."

            compile -library=libextras.a redboot_linux_exec.c
        }
    }
}
