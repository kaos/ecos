# ====================================================================
#
#      net_autotest.cdl
#
#      Networking autotest subsystem configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      hmt
# Original data:  hmt
# Contributors:
# Date:           2000-10-19
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_NET_AUTOTEST {
    display       "Networking autotest"
    doc           doc/index.html
    include_dir   net/autotest
    requires      CYGPKG_IO
    requires      CYGPKG_ISOINFRA
    requires      CYGPKG_LIBC_TIME
    requires      CYGPKG_ERROR
    requires      CYGPKG_MEMALLOC
    requires      CYGPKG_NET
    description   "Networking autotest facilities"

#    compile *NONE*

    cdl_option CYGPKG_NET_AUTOTEST_TESTS {
	display "Networking tests"
	flavor  data
	no_define
	calculated { "\
		tests/floodping.c \
		tests/floodpingmux.c \
		tests/route_3.c \
		tests/route_3_4.c \
		tests/route_4.c \
		tests/route_none.c \
		tests/slowping.c \
		tests/slowpingmux.c \
		tests/snmpwalk.c \
		tests/snmpmulti.c \
		tests/snmppings.c \
		tests/tftp_serv_get.c \
		tests/tftp_serv_put.c \
		tests/tftp_serv_g0.c \
		tests/tftp_serv_p0.c \
		tests/tftp_serv_g512.c \
		tests/tftp_serv_p512.c \
		tests/tftp_serv_g1M.c \
		tests/tftp_serv_p1M.c"
        }
	description   "
	This option specifies the set of tests
	for the networking package."
    }
	
    cdl_component CYGPKG_NET_AUTOTEST_OPTIONS {
        display "Networking support build options"
        flavor  none
	no_define

        cdl_option CYGPKG_NET_AUTOTEST_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building the autotest package.
	        These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_NET_AUTOTEST_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the autotest package. These flags are removed from
                the set of global flags if present."
        }
    }
}
