# ====================================================================
#
#      i386_pc_wallclock_drivers.cdl
#
#      Wallclock drivers - support for DS12887 RTC on the PC
#
# ====================================================================
#####COPYRIGHTBEGIN####
#
# -------------------------------------------
# The contents of this file are subject to the Red Hat eCos Public License
# Version 1.1 (the "License"); you may not use this file except in
# compliance with the License.  You may obtain a copy of the License at
# http://www.redhat.com/
#
# Software distributed under the License is distributed on an "AS IS"
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the
# License for the specific language governing rights and limitations under
# the License.
#
# The Original Code is eCos - Embedded Configurable Operating System,
# released September 30, 1998.
#
# The Initial Developer of the Original Code is Red Hat.
# Portions created by Red Hat are
# Copyright (C) 1998, 1999, 2000, 2001 Red Hat, Inc.
# All Rights Reserved.
# -------------------------------------------
#
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      rajt
# Contributors:   rajt
# Date:           2001-07-19
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVICES_WALLCLOCK_I386_PC {
    display       "PC board RTC Driver"
    description   "RTC driver for PC."

    parent        CYGPKG_IO_WALLCLOCK
    active_if   CYGPKG_IO_WALLCLOCK
    active_if     CYGPKG_HAL_I386_PC
    requires      CYGPKG_DEVICES_WALLCLOCK_DALLAS_DS12887

    include_dir   cyg/io

    define_proc {
        puts $::cdl_system_header "/***** PC RTC driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_DEVS_WALLCLOCK_DALLAS_12887_INL <cyg/io/devices_wallclock_i386_pc.inl>"
        puts $::cdl_system_header "#define CYGDAT_DEVS_WALLCLOCK_i386_PC_CFG <pkgconf/devices_wallclock_i386_pc.h>"
        puts $::cdl_system_header "/***** PC RTC driver proc output end  *****/"
    }

    cdl_option CYGDAT_DEVS_WALLCLOCK_I386_PC_RTC_ADDRESS_PORT {
    display         "IO port address of the ADDRESS register"
    flavor          data
        default_value 0x70
        description   "
              This option sets the io address of the address port for
              accessing the PC RTC"
    }

    cdl_option CYGDAT_DEVS_WALLCLOCK_I386_PC_RTC_DATA_PORT {
    display         "IO port address of the DATA register"
    flavor          data
        default_value 0x71
        description   "
              This option sets the io address of the data port for
              accessing the PC RTC"
    }
}
