# ====================================================================
#
#      io.cdl
#
#      eCos IO configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  gthomas
# Contributors:
# Date:           1999-07-07
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_IO {
    display       "I/O sub-system"
    doc           redirect/ecos-device-drivers.html
    include_dir   cyg/io
    requires      CYGPKG_ERROR
    description   "
        The eCos system is supplied with a number of different
        device drivers.  This option enables the basic I/O system
        support which is the basis for all drivers."

    compile       -library=libextras.a iosys.c ioinit.cxx io_diag.c
    compile       io_file.c

 
    cdl_option CYGDBG_IO_INIT {
        display       "Debug I/O sub-system"
        default_value 0
        description   "
            This option enables verbose messages to be displayed on the
            system 'diag' device during I/O system initialization."
   }

    cdl_option CYGPKG_IO_NFILE {
        display "Number of open files"
        flavor  data
        default_value 16
        description   "
            This option controls the number of open files."
    }
}
