# ====================================================================
#
#	ebsa285_eth_drivers.cdl
#
#	Ethernet drivers
#	Intel EBSA285 and PRO/100+ platform specific support
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      hmt
# Original data:  hmt
# Contributors:	  gthomas
# Date:           2000-02-01
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_ARM_EBSA285 {
    display       "Intel EBSA285 with PRO/100+ ethernet driver"

    parent        CYGPKG_NET_ETH_DRIVERS
    active_if     CYGPKG_NET_ETH_DRIVERS
    active_if     CYGPKG_HAL_ARM_EBSA285

    implements    CYGHWR_NET_DRIVER_ETH0
    implements    CYGHWR_NET_DRIVER_ETH1
    # yes, there should be two of these "implement"s
    implements    CYGHWR_NET_DRIVERS
    implements    CYGHWR_NET_DRIVERS
    include_dir   .
#    include_files ; # none _exported_ whatsoever
    description   "Ethernet driver for Intel EBSA285 with PRO/100+ boards."
    compile       -library=libextras.a if_ebsa285.c

    cdl_component CYGPKG_DEVS_ETH_ARM_EBSA285_OPTIONS {
        display "Intel EBSA285 with PRO/100+ ethernet driver build options"
        flavor  none
	no_define

        cdl_option CYGPKG_DEVS_ETH_ARM_EBSA285_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building the Intel EBSA285 with PRO/100+ ethernet driver
                package. These flags are used in addition to the set of
                global flags."
        }
    }
}

# EOF ebsa285_eth_drivers.cdl
