# ====================================================================
#
#      wallclock_stm32.cdl
#
#      Hardware support for STM32 on-chip RTC.
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2008 Free Software Foundation, Inc.                        
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Simon Kallweit
# Contributors:   
# Date:           2008-10-27
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_WALLCLOCK_STM32 {
    display       "STM32 RTC wallclock support"
    description   "
        Wallclock support for on-chip RTC on STM32 devices.driver for the
        STM32 controller and compatibles"

    parent        CYGPKG_IO_WALLCLOCK
    active_if     CYGPKG_IO_WALLCLOCK
    active_if     CYGPKG_HAL_CORTEXM_STM32

    compile       stm32_wallclock.cxx

    implements    CYGINT_WALLCLOCK_HW_IMPLEMENTATIONS
    active_if     CYGIMP_WALLCLOCK_HARDWARE
    implements    CYGINT_WALLCLOCK_SET_GET_MODE_SUPPORTED
    
    cdl_option CYGIMP_WALLCLOCK_HARDWARE {
        parent          CYGPKG_IO_WALLCLOCK_IMPLEMENTATION
        display         "Hardware wallclock"
        default_value   1
        implements      CYGINT_WALLCLOCK_IMPLEMENTATIONS
    }
    
    cdl_option CYGHWR_DEVS_WALLCLOCK_STM32_RTC_SOURCE {
        display             "RTC clock source"
        flavor              data
        default_value       { "LSE" }
        legal_values        { "LSE" "LSI" "HSE_128" }
    }
}
