# ====================================================================
#
#      hal_arm_arm9_innovator.cdl
#
#      TI Innovator platform HAL package configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Patrick Doyle <wpd@delcomsys.com>
# Contributors:   Patrick Doyle <wpd@delcomsys.com>
# Date:           2002-11-22
#
#####DESCRIPTIONEND####
#
# ====================================================================
cdl_package CYGPKG_HAL_ARM_ARM9_INNOVATOR {
    display       "Innovator"
    parent        CYGPKG_HAL_ARM_ARM9
    requires      CYGPKG_HAL_ARM_ARM9_ARM925T
    hardware
    include_dir   cyg/hal
    define_header hal_arm_arm9_innovator.h
    description   "
        This HAL platform package provides generic
        support for the OMAP Innovator platform."

    compile       innovator_misc.c hal_diag.c

    implements    CYGINT_HAL_DEBUG_GDB_STUBS
    implements    CYGINT_HAL_DEBUG_GDB_STUBS_BREAK
    implements    CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H   <pkgconf/hal_arm.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_VARIANT_H  <pkgconf/hal_arm_arm9.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_arm_arm9_innovator.h>"
	puts $::cdl_header "#define HAL_PLATFORM_CPU    \"ARM9\""
        puts $::cdl_header "#define HAL_PLATFORM_BOARD  \"Innovator\""
        puts $::cdl_header "#define HAL_PLATFORM_EXTRA  \"\""
        puts $::cdl_header "#define HAL_ARCH_PROGRAM_NEW_STACK innovator_program_new_stack"
        puts $::cdl_header "#define HAL_PLATFORM_MACHINE_TYPE  234"

    }

    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        default_value {"RAM"}
        legal_values  {"RAM" "ROM" }
	no_define
	define -file system.h CYG_HAL_STARTUP
        description   "
           When targetting the Innovator it is possible to build
           the system for either RAM bootstrap or ROM bootstrap(s). Select
           'RAM' when building programs to load into RAM using RedBoot.
           Select 'ROM' when building a stand-alone application
           which will be put into ROM, or for the special cases of
           building the eCos GDB stubs or RedBoot."

        cdl_option CYGPRI_HAL_ROM_MLT {
            display       "Memory Layout for ROM Startup"
            flavor        data
            legal_values  {"FLASH" "SRAM"}
            default_value {"FLASH"}
            description   "
                This option selects which memory layout file should be
		used when configuring the Innovator for ROM startup.
		The FLASH option selects the memory layout for an image
		stored at the beginning of the FLASH.  It should be
		used almost all of the time.

		The SRAM option is used to place the ROM image in
		internal SRAM.  It may be used in order to test startup
		code without burning the code into FLASH first." }
    }

    # Both PLLs are in bypass mode on startup.
    # FIXME: Add proper configury
    cdl_option CYGNUM_HAL_ARM_INNOVATOR_CPU_CLOCK {
        display       "CPU bus speed"
        flavor        data
        calculated    { 60000000 }
        description   "
            This is the actual CPU operating frequency.  Someday you
	    might be able to change this here."
    }

#    cdl_option CYGNUM_HAL_ARM_INNOVATOR_PERIPHERAL_CLOCK {
#        display       "Peripheral bus speed"
#        flavor        data
#        calculated    { CYGNUM_HAL_ARM_INNOVATOR_CPU_CLOCK / 2 }
#        description   "
#            This is the peripheral bus operating frequency
#	    (Traffic Controller)."
#    }
#
#    cdl_option CYGNUM_HAL_ARM_INNOVATOR_TIMER_PRESCALE {
#        display       "Timer prescale"
#        flavor        data
#        legal_values  0 to 255
#        default_value 16
#        description   "
#            This is the prescale value used on the clock used to drive
#            the kernel counter. Note that some parts of the code may fail
#            if this is changed due to over/underflows of expressions."
#    }
#
#    # Real-time clock/counter specifics
#    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
#        display       "Real-time clock constants.  WARNING -- the Real Time Clock is not fully supported (if at all) yet."
#        flavor        none
#        no_define
#    
#        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
#            display       "Real-time clock numerator"
#            flavor        data
#            calculated    1000000000
#        }
#        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
#            display       "Real-time clock denominator"
#            flavor        data
#            calculated    100
#        }
#        cdl_option CYGNUM_HAL_RTC_PERIOD {
#            display       "Real-time clock period"
#            flavor        data
#	    calculated	  1
##            calculated    (CYGNUM_HAL_ARM_INNOVATOR_PERIPHERAL_CLOCK/(CYGNUM_HAL_ARM_INNOVATOR_TIMER_PRESCALE*CYGNUM_HAL_RTC_DENOMINATOR))-1
#        }
#    }
#
#    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD {
#        display       "Diagnostic serial port baud rate"
#        flavor        data
#        legal_values  9600 19200 38400 57600 115200
#        default_value 115200
#        description   "
#            This option selects the baud rate used for the diagnostic port.
#            Note: this should match the value chosen for the GDB port if the
#            diagnostic and GDB port are the same."
#    }
#
#    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_BAUD {
#        display       "GDB serial port baud rate"
#        flavor        data
#        legal_values  9600 19200 38400 57600 115200
#        default_value 115200
#        description   "
#            This option selects the baud rate used for the diagnostic port.
#            Note: this should match the value chosen for the GDB port if the
#            diagnostic and GDB port are the same."
#    }
#
    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
        display      "Number of communication channels on the board"
        flavor       data
        calculated   1
    }
 
    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
        display          "Debug serial port"
        active_if        CYGPRI_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_CONFIGURABLE
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
            The Innovator has two serial ports.  When we add support
	    for the second one, you will be able to choose which one is
	    used to connect to a host running GDB."
     }

     cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_DEFAULT {
         display      "Default console channel."
         flavor       data
         legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
         calculated   0
     }
 
     cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
         display          "Diagnostic serial port"
         active_if        CYGPRI_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_CONFIGURABLE
         flavor data
         legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
         default_value    CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_DEFAULT
         description      "
            The Innovator has two serial ports.  When we add support
	    for the second one, you will be able to choose which one is
	    used for diagnostic output."
     }
 
    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        no_define
        description   "
	    Global build options including control over
	    compiler flags, linker flags and choice of toolchain."


        parent  CYGPKG_NONE

        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "arm-eabi"}
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { "-mcpu=arm9 -Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority" }
            description   "
                This option controls the global compiler flags which are used to
                compile all packages by default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { "--no-target-default-spec -Wl,--gc-sections -Wl,-static -g -O2 -nostdlib" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }

        cdl_option CYGBLD_BUILD_GDB_STUBS {
            display "Build GDB stub ROM image"
            default_value 0
            requires { CYG_HAL_STARTUP == "ROM" }
            requires CYGSEM_HAL_ROM_MONITOR
            requires CYGBLD_BUILD_COMMON_GDB_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT
            requires CYGDBG_HAL_DEBUG_GDB_THREAD_SUPPORT
            requires ! CYGDBG_HAL_COMMON_INTERRUPTS_SAVE_MINIMUM_CONTEXT
            requires ! CYGDBG_HAL_COMMON_CONTEXT_SAVE_MINIMUM
            no_define
            description "
                This option enables the building of the GDB stubs for the
                board. The common HAL controls takes care of most of the
                build process, but the final conversion from ELF image to
                binary data is handled by the platform CDL, allowing
                relocation of the data if necessary."

            make -priority 320 {
                <PREFIX>/bin/gdb_module.srec : <PREFIX>/bin/gdb_module.img
                $(OBJCOPY) --remove-section=.fixed_vectors $< gdb_module.tmp
            }
        }
    }

    cdl_component CYGPKG_HAL_ARM_ARM9_INNOVATOR_OPTIONS {
        display "Innovator build options"
        flavor  none
        no_define
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_HAL_ARM_ARM9_INNOVATOR_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the Innovator HAL. These flags are
		used in addition to the set of global flags."
        }

        cdl_option CYGPKG_HAL_ARM_ARM9_INNOVATOR_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the Innovator HAL. These flags are
		removed from the set of global flags if present."
        }

        cdl_option CYGPKG_HAL_ARM_ARM9_INNOVATOR_TESTS {
            display "Innovator tests"
            flavor  data
            no_define
            calculated { "" }
            description   "
                This option specifies the set of tests for the Innovator."
        }
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { CYG_HAL_STARTUP == "RAM" ? "arm_arm9_innovator_ram" : \
	                                        "arm_arm9_innovator_rom" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_arm9_innovator_ram.ldi>" : \
                         CYGPRI_HAL_ROM_MLT == "FLASH" ? "<pkgconf/mlt_arm_arm9_innovator_rom.ldi>" : \
                                                         "<pkgconf/mlt_arm_arm9_innovator_sram.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_arm9_innovator_ram.h>" : \
                         CYGPRI_HAL_ROM_MLT == "FLASH" ? "<pkgconf/mlt_arm_arm9_innovator_rom.h>" : \
                                                         "<pkgconf/mlt_arm_arm9_innovator_sram.h>" }
        }
    }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "ROM" }
        description   "
            Enable this option if this program is to be used as a ROM monitor,
            i.e. applications will be loaded into RAM on the board, and this
            ROM monitor may process exceptions or interrupts generated from the
            application. This enables features such as utilizing a separate
            interrupt stack when exceptions are generated."
    }

    cdl_option CYGSEM_HAL_USE_ROM_MONITOR {
         display       "Work with a ROM monitor"
         flavor        booldata
         legal_values  { "GDB_stubs" }
         default_value { CYG_HAL_STARTUP == "RAM" ? "GDB_stubs" : 0 }
         parent        CYGPKG_HAL_ROM_MONITOR
         requires      { CYG_HAL_STARTUP == "RAM" }
         description   "
             Support can be enabled for different varieties of ROM monitor.
             This support changes various eCos semantics such as the encoding
             of diagnostic output, or the overriding of hardware interrupt
             vectors.
             \"GDB_stubs\" provides support when GDB stubs are included in
             the ROM monitor or boot ROM."
     }

    cdl_component CYGPKG_REDBOOT_HAL_OPTIONS {
        display       "Redboot HAL options"
        flavor        none
        no_define
        parent        CYGPKG_REDBOOT
        active_if     CYGPKG_REDBOOT
        description   "
            This option lists the target's requirements for a valid Redboot
            configuration."

        # RedBoot details
        requires { CYGHWR_REDBOOT_ARM_LINUX_EXEC_ADDRESS_DEFAULT == 0x10008000 }
        define_proc {
            puts $::cdl_header "#define CYGHWR_REDBOOT_ARM_TRAMPOLINE_ADDRESS 0x00001f00"
        }

        cdl_option CYGBLD_BUILD_REDBOOT_BIN {
            display       "Build Redboot ROM binary image"
            active_if     CYGBLD_BUILD_REDBOOT
            default_value 1
            no_define
            description "This option enables the conversion of the Redboot ELF
                         image to the various relocated SREC images needed
                         for flash updating."

            compile -library=libextras.a redboot_cmds.c

            make -priority 325 {
                <PREFIX>/bin/redboot.bin : <PREFIX>/bin/redboot.elf
                $(OBJCOPY) --strip-debug $< $(@:.bin=.img) 
                $(OBJCOPY) -O srec $< $(@:.bin=.srec)
                $(OBJCOPY) -O binary $< $@
            }
        }
    }

}
