# ====================================================================
#
#      ser_sh_cq7708.cdl
#
#      eCos serial SH/CQ7708 configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Contributors:
# Date:           1999-07-08
#
#####DESCRIPTIONEND####
#
# ====================================================================


cdl_package CYGPKG_IO_SERIAL_SH_CQ7708 {
    display       "SH3 cq7708 serial device drivers"

    parent        CYGPKG_IO_SERIAL_DEVICES
    active_if     CYGPKG_IO_SERIAL
    active_if     CYGPKG_HAL_SH_SH7708_CQ7708

    requires      CYGPKG_ERROR
    include_dir   cyg/io

    description   "
           This option enables the serial device drivers for the
           CQ SH3 cq7708 board, based on the generic SH SCI driver."
    doc           redirect/ecos-device-drivers.html


    # FIXME: This really belongs in the SH_SCI package
    cdl_interface CYGINT_IO_SERIAL_SH_SCI_REQUIRED {
        display   "SH SCI driver required"
    }

    define_proc {
        puts $::cdl_system_header "/***** serial driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_SH_SCI_INL <cyg/io/sh_sh3_cq7708_sci.inl>"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_SH_SCI_CFG <pkgconf/io_serial_sh_cq7708.h>"
        puts $::cdl_system_header "/*****  serial driver proc output end  *****/"
    }

    cdl_component CYGPKG_IO_SERIAL_SH_CQ7708_SERIAL1 {
        display       "SH3 CQ7708 serial 1 device driver (SCI)"
        flavor        bool
        default_value 1
        description   "
            This option includes the serial device driver for the SCI
            port."

        implements CYGINT_IO_SERIAL_SH_SCI_REQUIRED

        cdl_option CYGDAT_IO_SERIAL_SH_CQ7708_SERIAL1_NAME {
            display       "Device name for SH3 CQ7708 SCI"
            flavor        data
            default_value {"\"/dev/ser1\""}
            description   "
                This option specifies the device name for the SCI port."
        }

        cdl_option CYGNUM_IO_SERIAL_SH_CQ7708_SERIAL1_BAUD {
            display       "Baud rate for the SH SCI driver"
            flavor        data
            legal_values  { 4800 9600 14400 19200 38400 57600 115200 }
            default_value 38400
            description   "
                This option specifies the default baud rate (speed)
                for the SCI port."
        }

        cdl_option CYGNUM_IO_SERIAL_SH_CQ7708_SERIAL1_BUFSIZE {
            display       "Buffer size for the SH SCI driver"
            flavor        data
            legal_values  0 to 8192
            default_value 128
            description   "
                This option specifies the size of the internal buffers
                used for the SCI port."
        }
    }

    cdl_component CYGPKG_IO_SERIAL_SH_CQ7708_TESTING {
        display    "Testing parameters"
        flavor     bool
        calculated 1
        no_define
        active_if  CYGPKG_IO_SERIAL_SH_CQ7708_SERIAL1

        define_proc {
            puts $::cdl_header "#define CYGPRI_SER_TEST_CRASH_ID \"sh-cq7708\""
            puts $::cdl_header "#define CYGPRI_SER_TEST_SER_DEV  CYGDAT_IO_SERIAL_SH_CQ7708_SERIAL1_NAME"
            puts $::cdl_header "#define CYGPRI_SER_TEST_TTY_DEV  \"/dev/tty1\""
        }
    }
}
# EOF ser_sh_cq7708.cdl
