# ====================================================================
#
#      hal.cdl
#
#      HAL configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      bartv
# Original data:  nickg,jskov,jlarmour
# Contributors:
# Date:           1999-06-13
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL {
    display       "eCos HAL"
    include_dir   cyg/hal
    description   "
        The eCos HAL package provide a porting layer for
        higher-level parts of the system such as the kernel and the
        C library. Each installation should have HAL packages for
        one or more architectures, and for each architecture there
        may be one or more supported platforms. It is necessary to
        select one target architecture and one platform for that
        architecture. There are also a number of configuration
        options that are common to all HAL packages."
    doc           redirect/the-ecos-hardware-abstraction-layer-hal.html

    compile       generic-stub.c thread-packets.c hal_stub.c drv_api.c
    compile       -library=libextras.a dummy.c

    make -priority 250 {
        <PREFIX>/lib/extras.o: <PREFIX>/lib/libextras.a
        $(CC) $(CFLAGS) -nostdlib -Wl,-r -Wl,--whole-archive -o $@ $<
    }   


    cdl_component CYGPKG_HAL_COMMON {
        display       "Platform-independent HAL options"
        flavor        none
        description   "
            A number of configuration options are common to most or all
            HAL packages, for example options controlling how much state
            should be saved during a context switch. The implementations
            of these options will vary from architecture to architecture."

        script        common.cdl
    }

    cdl_component CYGPKG_HAL_COMMON_INTERRUPTS {
        display       "HAL interrupt handling"
        flavor        none
        description   "
            A number of configuration options related to interrupt
            handling are common to most or all HAL packages, even though
            the implementations will vary from architecture to
            architecture."

        script        interrupts.cdl
    }

    cdl_component CYGPKG_HAL_COMMON_CONTEXT {
        display       "HAL context switch support"
        flavor        none
        description   "
            A number of configuration options related to thread contexts
            are common to most or all HAL packages, even though the
            implementations will vary from architecture to architecture."

        cdl_option CYGDBG_HAL_COMMON_CONTEXT_SAVE_MINIMUM {
            display       "Use minimum thread context"
            parent        CYGPKG_HAL_COMMON_CONTEXT
            default_value 1
            description   "
                The thread context switch code can exploit the calling
                conventions defined for a given architecture to reduce the
                amount of state that has to be saved during a context
                switch. Generally this improves performance and reduces
                code size. However it can make source-level debugging more
                difficult."
        }
    }

    cdl_component CYGPKG_HAL_DEBUG {
        display       "Source-level debugging support"
        flavor        none
        description   "
            If the source level debugger gdb is to be used for debugging
            application code then it may be necessary to configure in support
            for this in the HAL."

        script        debugging.cdl
    }

    cdl_component CYGPKG_HAL_ROM_MONITOR {
        display       "ROM monitor support"
        flavor        none
        no_define
        description   "
            Support for ROM monitors can be built in to your application. 
            It may also be relevant to build your application as a ROM monitor
            itself. Such options are contained here if relevant for your chosen
            platform. The options and ROM monitors available to choose are
            platform-dependent."


        cdl_option CYGBLD_BUILD_COMMON_GDB_STUBS {
            display "Build common GDB stub ROM image"
            default_value 0
            parent  CYGBLD_GLOBAL_OPTIONS
            requires CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
            no_define
            description "
                Unless a target board has specific requirements to the
                stub implementation, it can use a simple common stub.
                This option, which gets enabled by platform HALs as
                appropriate, controls the building of the common stub."
                         
            make -priority 315 {
                <PREFIX>/bin/gdb_module.img : <PACKAGE>/src/stubrom/stubrom.c <PREFIX>/lib/extras.o <PREFIX>/lib/libtarget.a <PREFIX>/lib/target.ld <PREFIX>/lib/vectors.o
                @sh -c "mkdir -p src/stubrom $(dir $@)"
                $(CC) -c $(INCLUDE_PATH) -Wp,-MD,deps.tmp -I$(dir $<) $(CFLAGS) -o src/stubrom/gdb_module.o $<
                @echo $@ ": \\" > $(notdir $@).deps
                @echo $(wildcard $(PREFIX)/lib/*) " \\" >> $(notdir $@).deps
                @tail +2 deps.tmp >> $(notdir $@).deps
                @echo >> $(notdir $@).deps
                @rm deps.tmp
                $(CC) $(LDFLAGS) -L$(PREFIX)/lib -Ttarget.ld -o $@ src/stubrom/gdb_module.o
            }
        }


    }

    define_proc {
        puts $::cdl_header "/***** proc output start *****/"
        puts $::cdl_header "#include <pkgconf/system.h>"

        puts $::cdl_header "#include CYGBLD_HAL_TARGET_H"
        puts $::cdl_header "#include CYGBLD_HAL_PLATFORM_H"

        puts $::cdl_header "/****** proc output end ******/"

    }

    cdl_option CYGPKG_HAL_TESTS {
        display "Common HAL tests"
        flavor  data
        no_define
        calculated { "tests/cache tests/context tests/intr" }
        description   "
            This option specifies the set of tests for the common HAL."
    }
}
