# ====================================================================
#
#      hal_arm_sa11x0.cdl
#
#      ARM SA11x0 architectural HAL package configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Original data:  gthomas
# Contributors:
# Date:           2000-05-08
#
#####DESCRIPTIONEND####
#
# ====================================================================
cdl_package CYGPKG_HAL_ARM_SA11X0 {
    display       "ARM SA11X0 architecture"
    parent        CYGPKG_HAL_ARM
    hardware
    include_dir   cyg/hal
    define_header hal_arm_sa11x0.h
    description   "
        This HAL variant package provides generic
        support for the Intel StrongARM SA11x0 processors. It is also
        necessary to select a specific target platform HAL
        package."


    compile       hal_diag.c sa11x0_misc.c

    cdl_option CYGHWR_HAL_ARM_SA11X0_PROCESSOR_CLOCK {
        display       "Processor clock rate"
        flavor        data
        legal_values  59000 73700 88500 103200 118000 132700 147500 162200 176900 191700 206400 221200
        default_value 221200
        description   "
           The SA-1100 processor can run at various frequencies.
           These values are expressed in KHz.  Note that there are
           several steppings of the SA-1100 rated to run at different
           maximum frequencies.  Check the specs to make sure that your
           particular processor can run at the rate you select here."
    }

    # Real-time clock/counter specifics
    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants"
        flavor        none
        no_define
    
        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            calculated    1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            calculated    100
        }
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
            calculated    36864        ;# Clock for OS Timer is 3.6864MHz
        }
    }

}
