# ====================================================================
#
#      net.cdl
#
#      Networking configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000, 2001 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Original data:  gthomas
# Contributors:
# Date:           1999-11-29
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_NET {
    display       "Networking"
    doc           doc/index.html
    include_dir   .
    requires      CYGPKG_IO
    requires      CYGPKG_ISOINFRA
    requires      CYGINT_ISO_C_TIME_TYPES
    requires      CYGINT_ISO_STRERROR
    requires      CYGINT_ISO_ERRNO
    requires      CYGINT_ISO_ERRNO_CODES
    requires      CYGINT_ISO_MALLOC
    description   "Basic networking support, including TCP/IP."

    cdl_interface     CYGPKG_NET_DRIVER_FRAMEWORK {
        display   "Suitable driver framework interface, used by network package"
        description "
          In order to decouple the network stack from driver specifics, the
          driver framework must be defined in a separate package."
    }

    # Export our types to <sys/types.h>
    implements    CYGINT_ISO_BSDTYPES
    requires      { CYGBLD_ISO_BSDTYPES_HEADER == "<sys/bsdtypes.h>" }
    implements    CYGINT_ISO_NETDB_PROTO
    implements    CYGINT_ISO_NETDB_SERV
    requires      { CYGBLD_ISO_NETDB_PROTO_HEADER == "<net/netdb.h>" }
    requires      { CYGBLD_ISO_NETDB_SERV_HEADER == "<net/netdb.h>" }
    
    compile ecos/support.c \
        ecos/synch.c \
        ecos/timeout.c \
        ecos/init.cxx \
        sys/kern/uipc_mbuf.c \
        sys/kern/uipc_domain.c \
        sys/kern/uipc_socket.c \
        sys/kern/uipc_socket2.c \
        sys/kern/kern_subr.c \
        sys/net/if.c \
        sys/net/rtsock.c \
        sys/net/raw_cb.c \
        sys/net/raw_usrreq.c \
        sys/net/route.c \
        sys/net/radix.c \
        sys/net/if_ethersubr.c \
        sys/net/if_loop.c \
        sys/netinet/igmp.c \
        sys/netinet/raw_ip.c \
        sys/netinet/in.c  \
        sys/netinet/in_cksum.c \
        sys/netinet/in_pcb.c \
        sys/netinet/in_proto.c \
        sys/netinet/ip_id.c \
        sys/netinet/ip_icmp.c \
        sys/netinet/ip_input.c \
        sys/netinet/ip_output.c \
        sys/netinet/if_ether.c \
        sys/netinet/udp_usrreq.c \
        sys/netinet/tcp_input.c \
        sys/netinet/tcp_output.c \
        sys/netinet/tcp_subr.c \
        sys/netinet/tcp_debug.c \
        sys/netinet/tcp_usrreq.c \
        sys/netinet/tcp_timer.c \
        lib/inet_addr.c \
        lib/bootp_support.c \
        lib/dhcp_support.c \
        lib/dhcp_prot.c \
        lib/network_support.c \
        lib/getproto.c \
        lib/getserv.c

    cdl_option CYGPKG_NET_API_LOCAL {
        display "Implement the socket API locally"
        flavor bool
        active_if !CYGPKG_IO_FILEIO
        default_value 1
        implements CYGINT_ISO_SELECT
        
        compile sys/kern/uipc_syscalls.c \
        sys/kern/sys_socket.c \
        sys/kern/sys_generic.c \
        lib/socket.c \
        lib/close.c \
        lib/read.c \
        lib/write.c \
        lib/bind.c \
        lib/connect.c \
        lib/accept.c \
        lib/listen.c \
        lib/shutdown.c \
        lib/sendto.c \
        lib/recvfrom.c \
        lib/getsockname.c \
        lib/getpeername.c \
        lib/getsockopt.c \
        lib/setsockopt.c \
        lib/ioctl.c \
        lib/select.c

        description "
            This option controls support for the network-stack supplied
            API."
    }

    cdl_option CYGPKG_NET_API_FILEIO {
        display "Implement the socket API via Fileio package"
        active_if CYGPKG_IO_FILEIO
        default_value 1

        compile -library=libextras.a sys/kern/sockio.c

        description "
            This option controls support for the fileio subsystem supplied API."
    }

    cdl_component CYGPKG_NET_INET {
        display "INET support"
        flavor  bool
        no_define
        default_value 1
        description   "
            This option enables support for INET (IP) network processing."
        define INET

        cdl_option CYGPKG_NET_INET6 {
            display "IPv6 support"
            flavor  bool
            default_value 0
            description   "
                This option enables support for new IPv6."
            define INET6
        }

        cdl_option CYGPKG_NET_ROUTING {
            display "Routing support"
            flavor  bool
            no_define
            default_value 0
            description   "
                This option enables support for packet routing."
            define MROUTING
        }

    }

    cdl_component CYGPKG_NET_TFTP {
        display        "TFTP (RFC-1350) support"
        flavor         bool
        default_value  1
        compile        lib/tftp_client.c \
                       lib/tftp_server.c
        description    "
          This option provides additional library support for
          the TFTP (Trivial File Transfer Protocol)."

        cdl_option CYGPKG_NET_TFTPD_THREAD_PRIORITY {
            display "Priority level for TFTP daemon thread."
            flavor  data
            default_value 10
            description   "
            This option allows the thread priority level used by the
            TFTP server thread to be adjusted by the user.  It should be set
            high enough that sufficient CPU resources are available to
            process network data, but may be adjusted so that application
            threads can have precedence over TFTP server processing."
        }

        cdl_option CYGPKG_NET_TFTP_FILE_ACCESS {
            display       "File I/O functions for TFTP server"
            flavor        bool
            default_value 1
            compile       lib/tftp_dummy_file.c
            description   "
              Minimal in-memory file I/O support for TFTP server."
        }
    }

    cdl_component CYGPKG_NET_DHCP {
        display "Use full DHCP instead of BOOTP"
        active_if (CYGHWR_NET_DRIVERS > 0)
        flavor bool
        default_value 1
        description "
            Provide DHCP for initializing the IP address
            of network interfaces.  The DHCP client is capable of falling
            back to BOOTP usage if the server does not support DHCP, so it
            should never be necessary to disable this option.  However,
            depending on other configuration the DHCP client may provide or
            require a kernel thread of its own; this consumes quite a lot
            of resource which a BOOTP solution does not require."

        cdl_option CYGOPT_NET_DHCP_DHCP_THREAD {
            display "DHCP management thread"
            flavor bool
            default_value 1
            description "
                Provide a separate thread to renew DHCP leases; otherwise
                the application MUST periodically examine the semaphore
                dhcp_needs_attention and call dhcp_bind() if it is
                signalled.  If enabled, this thread does all that for you.
                Independent of this option, initialization of the
                interfaces still occurs in init_all_network_interfaces()
                and your startup code must call that.  It will start the
                DHCP management thread if necessary.  If a lease fails to
                be renewed, the management thread will shut down all
                interfaces and attempt to initialize all the interfaces
                again from scratch.  This may cause application problems,
                in which case managing the DHCP state in an application
                aware thread is recommended.  See comments in dhcp.h"
        }

        cdl_option CYGOPT_NET_DHCP_DHCP_THREAD_PARAM {
            display "DHCP management thread loops forever"
            flavor  data
            default_value 1
            active_if CYGOPT_NET_DHCP_DHCP_THREAD
            description "
                If the parameter is nonzero, it loops forever; if zero,
                the thread exits if a lease expires, and the application
                must detect this and tidy up or reboot the whole machine."
        }
        cdl_option CYGPKG_NET_DHCP_THREAD_PRIORITY {
            display "DHCP management thread priority"
            flavor  data
            default_value CYGPKG_NET_THREAD_PRIORITY + 1
            active_if CYGOPT_NET_DHCP_DHCP_THREAD
            description "
            This option sets the thread priority level used by the DHCP
            management thread.  It should be high enough that it can run
            when necessary, but it does not need to be as high as the
            network thread itself."
        }
    }

#    cdl_option CYGPKG_NET_SYSCTL {
#        display "Support BSD 'sysctl()' function"
#        flavor  bool
#        default_value 0
#        description   "
#            This option includes support for the 'sysctl()' functions."
#    }

    cdl_option CYGPKG_NET_THREAD_PRIORITY {
        display "Priority level for backgound network processing."
        flavor  data
        default_value 7
        description   "
            This option allows the thread priority level used by the
        networking stack to be adjusted by the user.  It should be set
        high enough that sufficient CPU resources are available to
        process network data, but may be adjusted so that application
        threads can have precedence over network processing."
    }

    cdl_option CYGPKG_NET_FAST_THREAD_PRIORITY {
        display "Priority level for fast network processing."
        flavor  data
        default_value CYGPKG_NET_THREAD_PRIORITY - 1
        description   "
            This option sets the thread priority level used by the fast
        network thread.  The fast network thread runs often but briefly, to
        service network device interrupts and network timeout events.  This
        thread should have higher priority than the background network
        thread.  It is reasonable to set this thread's priority higher than
        application threads for best network throughput, or to set it lower
        than application threads for best latency for those application
        threads themselves, potentially at a cost to network throughput."
    }

    cdl_component CYGPKG_NET_FAST_THREAD_TICKLE_DEVS {
        display "Fast network processing thread 'tickles' drivers"
        default_value 1
        description "
            If this is enabled, the fast network thread will tickle the
            device(s) periodically, to unblock them when the hardware has
            become wedged due to a lost interrupt or other hardware
            race-condition type problem.
            This is not necessary if a networked app is running which sends
            packets itself often - or
            uses TCP, or any similar protocol which exchanges keep-alive
            packets periodically and often enough.
            Trying to send a packet passes control into the driver; this is
            sufficient to detect and unblock jammed hardware."

        cdl_option CYGNUM_NET_FAST_THREAD_TICKLE_DEVS_DELAY {
            display "Delay in kernel clocks of tickle loop"
            flavor data
            default_value 50
            description "
                The default is 50, which will usually mean a delay between
                tests for 'stuck' devices of 500mS, that is half a second.
	        The overhead only applies if no network activity occurred,
	        so it may be acceptable to make this value very small,
                where high CPU load does not matter during network idle
                periods, or very large if your application tries often to
                send packets itself."
        }
    }

    cdl_option CYGPKG_NET_NBPF {
        display "Number of BPF filters"
        flavor  data
        default_value 0
        description   "
            This option controls the number of active BPF filters."
        define NBPFILTER
    }

    cdl_component CYGPKG_NET_BRIDGE {
         display "Built-in ethernet bridge code"
         default_value 0
         implements CYGINT_NET_BRIDGE_HANDLER
     no_define
         description   "
             This option controls whether to include the built-in code for
             the Ethernet bridge."
     compile sys/net/if_bridge.c

         cdl_option CYGNUM_NET_BRIDGES {
             display "Number of Ethernet bridges"
             flavor  data
             default_value 1
             legal_values 1 to 999999
         }
    }

    cdl_interface CYGINT_NET_BRIDGE_HANDLER {
        display "Support for ethernet bridges in the IP stack"
        define NBRIDGE
            description "
              This interface controls whether calls to bridge code are made
              from the IP stack; these are needed if the built-in bridge code
              is used, but they can also be enabled in order to call different
              bridge code from an external component."
    }

    cdl_option CYGPKG_NET_NGIF {
        display "Number of GIF things"
        flavor  data
        default_value 0
        description   "
            This option controls the number of active GIF things."
        define NGIF
    }

    cdl_option CYGPKG_NET_NLOOP {
        display "Number of loopback interfaces"
        flavor  data
        default_value 1
        requires { (CYGPKG_NET_NLOOP > 1) ? CYGPKG_LIBC_STDIO : 1  }
        description   "
            This option controls the number of loopback, i.e. local, interfaces.
            There is seldom need for this value to be anything other than one.
            If a different value is required, then the C library STDIO package
            is required for sprintf()."
        define NLOOP
    }

    cdl_option CYGPKG_NET_MEM_USAGE {
        display "Memory designated for networking buffers."
        flavor  data
        default_value 256*1024
        description   "
            This option controls the amount of memory pre-allocated
        for buffers used by the networking code."
    }

    cdl_option CYGPKG_NET_NUM_WAKEUP_EVENTS {
        display "Number of supported pending network events"
        flavor  data
        default_value 8
        description   "
            This option controls the number of pending network events
        used by the networking code."
    }

    cdl_component CYGPKG_NET_DEBUG {
        display       "Debug output"
        default_value 0 
        description   "
                This component controls whether there is diagnostic output
                for stack operations. Options within this component allow
                even more verbose output for certain areas."

        cdl_option CYGDBG_NET_DHCP_CHATTER {
                display       "Extra debug output for DHCP"
                default_value 0
        }
    }

    cdl_component CYGPKG_NET_OPTIONS {
        display "Networking support build options"
        flavor  none
        no_define

        cdl_option CYGPKG_NET_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS -D__INSIDE_NET" }
            description   "
                This option modifies the set of compiler flags for
                building the networking package.
                These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_NET_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the networking package. These flags are removed from
                the set of global flags if present."
        }
    }

    cdl_component CYGPKG_NET_BUILD_TESTS {
        display "Build networking tests (demo programs)"
        flavor  bool
        no_define
        default_value 0
        description   "
        This option enables the building of additional network tests
        which at this time are just demos; otherwise only loopback
        interface tests will be built."

        cdl_option CYGPKG_NET_TESTS {
            display "Networking tests"
            flavor  data
            no_define
            calculated { CYGPKG_NET_BUILD_TESTS ? \
                    "tests/mbuf_test \
                    tests/socket_test \
                    tests/ftp_test \
                    tests/server_test \
                    tests/nc_test_slave \
                    tests/tftp_client_test \
                    tests/tftp_server_test \
                    tests/tcp_echo \
                    tests/set_mac_address \
                    tests/bridge \
                    tests/flood \
                    tests/ping_test \
                    tests/dhcp_test \
                    tests/ping_lo_test \
                    tests/tcp_lo_test \
                    tests/udp_lo_test \
                    tests/multi_lo_select \
                    tests/tcp_lo_select"
            :
                    "tests/ping_lo_test \
                    tests/tcp_lo_test \
                    tests/udp_lo_test \
                    tests/multi_lo_select \
                    tests/tcp_lo_select"
        }
            description   "
            This option specifies the set of tests
            for the networking package."
        }
        
        cdl_option CYGPKG_NET_TESTS_USE_RT_TEST_HARNESS {
            display "Use real-time response test harness (if available)"
            default_value 0
            description "
                    Platform and/or ethernet device driver packages may
                    provide a test harness to verify that interrupts are
                    not disabled or flooded for too long during a test.  If
                    such is provided, CYGTST_DEVS_ETH_TEST_NET_REALTIME is
                    defined and can be #include'd to acquire the support.
                    Some tests in the TCP/IP stack can use this harness;
                    this option controls whether they do.  The StrongARM
                    EBSA285 Ethernet device driver is one package that
                    provides such a harness.  See the file
                    tests/test_net_realtime.h in there for details."
        }
    }

# Description and control over different interfaces

    cdl_interface CYGHWR_NET_DRIVERS {
        display "Network drivers"
    }

    cdl_interface CYGHWR_NET_DRIVER_ETH0 {
        display "Does the hardware provide an 'eth0' device?"
        requires { CYGHWR_NET_DRIVER_ETH0 <= 1 }
        flavor   bool
    }

    cdl_component CYGHWR_NET_DRIVER_ETH0_SETUP_OPTIONS {
        display "Initialization options for 'eth0'"
        active_if (CYGHWR_NET_DRIVER_ETH0 == 1)
        flavor none
        no_define

        cdl_interface CYGHWR_NET_DRIVER_ETH0_SETUP {
            display "Initialization options for 'eth0'"
            requires 1 == CYGHWR_NET_DRIVER_ETH0_SETUP
            no_define
        }

        cdl_component CYGHWR_NET_DRIVER_ETH0_MANUAL {
            display "Initialize 'eth0' manually?"
            default_value 0
            implements CYGHWR_NET_DRIVER_ETH0_SETUP
            description "
                If this option is selected, the eCos library provides no
                initialization code for this interface; you must perform
                all the initialization in the application, by means of
                appropriate ioctl() calls, or by calling init_net() with an
                appropriate bootp record you have constructed yourself."
        }

        cdl_component CYGHWR_NET_DRIVER_ETH0_BOOTP {
            display "Use BOOTP/DHCP to initialize 'eth0'?"
            default_value 1
            implements CYGHWR_NET_DRIVER_ETH0_SETUP     
            description "
                If this option is selected, init_all_network_interfaces()
                will use DHCP or BOOTP to acquire initialization data for
                this interface, and then set it up accordingly."

            cdl_option CYGHWR_NET_DRIVER_ETH0_DHCP {
                display "Use DHCP rather than BOOTP for 'eth0'?"
                flavor  bool
                default_value 1
                active_if CYGPKG_NET_DHCP
            }

            cdl_option CYGHWR_NET_DRIVER_ETH0_BOOTP_SHOW {
                display "Show BOOTP/DHCP initialization values?"
                flavor  bool
                default_value 1
            }
        }

        cdl_component CYGHWR_NET_DRIVER_ETH0_ADDRS {
            display "Address setups for 'eth0'"
            implements CYGHWR_NET_DRIVER_ETH0_SETUP     
            no_define

            description "
                These options let you configure all the initialization data
                that init_all_network_interfaces() will use
                for 'eth0' statically.  Be careful when doing this, because
                if you run the same application image on multiple boards,
                they will have identical IP addresses and so on; this is a
                Bad Thing.
                The values you set are inserted in a bootp-style record
                that is fed into a common setup routine to configure the
                interface.  That routine does not in fact use the 'Server
                IP address' field.
                The bootp record is also available to application code, and
                some eCos networking test programs use the 'Server IP
                address' field to mean 'a machine we can interact with' for
                example to ping or perform ftp with.  That is the rationale
                for its inclusion here.
                The gateway address is used to set up a default route if
                nonzero.  If you have more than one interface, setting up
                more than one default route is will cause malfunctions.  A
                gateway address of 0.0.0.0 can be set to prevent that route
                setup.  Of course, your application can add real routes
                once the interface(s) initialization is complete."

            cdl_option CYGHWR_NET_DRIVER_ETH0_ADDRS_IP {
                display "IP address for 'eth0'"
                flavor  data
                default_value { "192.168.1.2" }
            }

            cdl_option CYGHWR_NET_DRIVER_ETH0_ADDRS_NETMASK {
                display "Network mask address for 'eth0'"
                flavor  data
                default_value { "255.255.255.0" }
            }

            cdl_option CYGHWR_NET_DRIVER_ETH0_ADDRS_BROADCAST {
                display "Broadcast address for 'eth0'"
                flavor  data
                default_value { "192.168.1.255" }
            }

            cdl_option CYGHWR_NET_DRIVER_ETH0_ADDRS_GATEWAY {
                display "Gateway/router IP address for 'eth0'"
                flavor  data
                default_value { "192.168.1.1" }
            }

            cdl_option CYGHWR_NET_DRIVER_ETH0_ADDRS_SERVER {
                display "Server IP address for 'eth0'"
                flavor  data
                default_value { "192.168.1.101" }
            }
        }
    }

    cdl_interface CYGHWR_NET_DRIVER_ETH1 {
        display "Does the hardware provide an 'eth1' device?"
        requires { CYGHWR_NET_DRIVER_ETH1 <= 1 }
        flavor   bool
    }

    cdl_component CYGHWR_NET_DRIVER_ETH1_SETUP_OPTIONS {
        display "Initialization options for 'eth1'"
        active_if (CYGHWR_NET_DRIVER_ETH1 == 1)
        flavor none
        no_define

        cdl_interface CYGHWR_NET_DRIVER_ETH1_SETUP {
            display "Initialization options for 'eth1'"
            requires 1 == CYGHWR_NET_DRIVER_ETH1_SETUP
            no_define
        }

        cdl_component CYGHWR_NET_DRIVER_ETH1_MANUAL {
            display "Initialize 'eth1' manually?"
            default_value 0
            implements CYGHWR_NET_DRIVER_ETH1_SETUP     
            description "
                If this option is selected, the eCos library provides no
                initialization code for this interface; you must perform
                all the initialization in the application, by means of
                appropriate ioctl() calls, or by calling init_net() with an
                appropriate bootp record you have constructed yourself."
        }

        cdl_component CYGHWR_NET_DRIVER_ETH1_BOOTP {
            display "Use BOOTP/DHCP to initialize 'eth1'?"
            default_value 1
            implements CYGHWR_NET_DRIVER_ETH1_SETUP     
            description "
                If this option is selected, init_all_network_interfaces()
                will use DHCP or BOOTP to acquire initialization data for
                this interface, and then set it up accordingly."

            cdl_option CYGHWR_NET_DRIVER_ETH1_DHCP {
                display "Use DHCP rather than BOOTP for 'eth1'?"
                flavor  bool
                default_value 1
                active_if CYGPKG_NET_DHCP
            }

            cdl_option CYGHWR_NET_DRIVER_ETH1_BOOTP_SHOW {
                display "Show BOOTP/DHCP initialization values?"
                flavor  bool
                default_value 1
            }
        }

        cdl_component CYGHWR_NET_DRIVER_ETH1_ADDRS {
            display "Address setups for 'eth1'"
            implements CYGHWR_NET_DRIVER_ETH1_SETUP     
            no_define

            description "
                These options let you configure all the initialization data
                that init_all_network_interfaces() will use
                for 'eth1' statically.  Be careful when doing this, because
                if you run the same application image on multiple boards,
                they will have identical IP addresses and so on; this is a
                Bad Thing.
                The values you set are inserted in a bootp-style record
                that is fed into a common setup routine to configure the
                interface.  That routine does not in fact use the 'Server
                IP address' field.
                The bootp record is also available to application code, and
                some eCos networking test programs use the 'Server IP
                address' field to mean 'a machine we can interact with' for
                example to ping or perform ftp with.  That is the rationale
                for its inclusion here.
                The gateway address is used to set up a default route if
                nonzero.  If you have more than one interface, setting up
                more than one default route is will cause malfunctions.  A
                gateway address of 0.0.0.0 can be set to prevent that route
                setup.  Of course, your application can add real routes
                once the interface(s) initialization is complete.
                This interface 'eth1' has no route set up in the default
                configuration."

            cdl_option CYGHWR_NET_DRIVER_ETH1_ADDRS_IP {
                display "IP address for 'eth1'"
                flavor  data
                default_value { "192.168.1.2" }
            }

            cdl_option CYGHWR_NET_DRIVER_ETH1_ADDRS_NETMASK {
                display "Network mask address for 'eth1'"
                flavor  data
                default_value { "255.255.255.0" }
            }

            cdl_option CYGHWR_NET_DRIVER_ETH1_ADDRS_BROADCAST {
                display "Broadcast address for 'eth1'"
                flavor  data
                default_value { "192.168.1.255" }
            }

            cdl_option CYGHWR_NET_DRIVER_ETH1_ADDRS_GATEWAY {
                display "Gateway/router IP address for 'eth1'"
                flavor  data
                default_value { "0.0.0.0" }
            }

            cdl_option CYGHWR_NET_DRIVER_ETH1_ADDRS_SERVER {
                display "Server IP address for 'eth1'"
                flavor  data
                default_value { "192.168.1.101" }
            }
        }
    }
}
