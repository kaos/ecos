# ====================================================================
#
#      posix.cdl
#
#      POSIX layer configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000, 2001 Red Hat, Inc.      
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      nickg
# Contributors:
# Date:           2000-3-28
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_POSIX {
    display        "POSIX compatibility layer"
    description    "This package enables the POSIX compatibility
                    layer that implements IEEE 1003.1."
    include_dir    cyg/posix
    
    requires       CYGPKG_KERNEL
    requires       CYGPKG_ISOINFRA
    requires       CYGPKG_ERROR
    requires       CYGINT_ISO_ERRNO
    requires       CYGINT_ISO_ERRNO_CODES
    requires       CYGIMP_KERNEL_SCHED_SORTED_QUEUES

    implements     CYGINT_ISO_SCHED_IMPL
    implements     CYGINT_ISO_POSIX_LIMITS
    requires       { CYGBLD_ISO_POSIX_LIMITS_HEADER == \
                         "<cyg/posix/limits.h>" }
    
    compile        mqueue.cxx mutex.cxx sem.cxx misc.cxx
    compile       -library=libextras.a startup.cxx

    # ----------------------------------------------------------------
    # Scheduling component
    
    cdl_component CYGPKG_POSIX_SCHED {
	display          "POSIX scheduling configuration"
	flavor           bool
	default_value    1
	description      "This component provides controls over scheduling
	                  in POSIX."
        requires         CYGPKG_POSIX_TIMERS
        compile          sched.cxx

	cdl_option _POSIX_PRIORITY_SCHEDULING {
	    display       "POSIX priority scheduling feature test macro"
	    flavor        bool
	    calculated    1
	    requires      CYGSEM_KERNEL_SCHED_MLQUEUE
	    description   "This option defines the POSIX feature test macro
	                   that indicates that priority scheduling is present.
	                   This should not be undefined."
	}
    }

    # ----------------------------------------------------------------
    # Pthreads component

    cdl_component CYGPKG_POSIX_PTHREAD {
	display          "POSIX pthread configuration"
	flavor           bool
	default_value    1
	description      "This component provides configuration controls for
	                  the POSIX pthreads package."
        compile          pthread.cxx
	script           pthread.cdl
    }

    # ----------------------------------------------------------------
    # Timers component

    cdl_option CYGPKG_POSIX_TIMERS {
	display          "POSIX timers"
	flavor           bool
	default_value    1
        implements       CYGINT_ISO_POSIX_TIMER_TYPES
        implements       CYGINT_ISO_POSIX_TIMERS
        implements       CYGINT_ISO_POSIX_TIMER_OPS
        requires         { CYGBLD_ISO_POSIX_TIMER_TYPES_HEADER == \
                             "<cyg/posix/time.h>" }
        requires         { CYGBLD_ISO_POSIX_TIMERS_HEADER == \
                             "<cyg/posix/time.h>" }
        requires         CYGPKG_KERNEL
        requires         CYGVAR_KERNEL_COUNTERS_CLOCK
        requires         CYGPKG_POSIX_PTHREAD
        compile          time.cxx
	description      "This component provides configuration controls for
	                  the POSIX timers."
    }

    # ----------------------------------------------------------------
    # Semaphores component

    cdl_option CYGPKG_POSIX_SEMAPHORES {
	display          "POSIX semaphores"
	flavor           bool
	default_value    1
        implements       CYGINT_ISO_SEMAPHORES
        requires         { CYGBLD_ISO_SEMAPHORES_HEADER == \
                             "<cyg/posix/semaphore.h>" }
	description      "This component provides configuration controls for
	                  POSIX semaphores."
    }

    # ----------------------------------------------------------------
    # Message queues component

    cdl_component CYGPKG_POSIX_MQUEUES {
	display          "POSIX message queues"
	flavor           bool
	default_value    1
        implements       CYGINT_ISO_MQUEUE
        requires         CYGPKG_KERNEL
        requires         CYGINT_ISO_MALLOC
        requires         CYGINT_ISO_ERRNO
        requires         CYGINT_ISO_STRING_STRFUNCS
	description      "This component provides configuration controls for
	                  POSIX message queues."

        cdl_option CYGNUM_POSIX_MQUEUE_OPEN_MAX {
            display          "Maximum number of message queues"
            flavor           data
            default_value    8
            legal_values     1 to 999999
        }

        cdl_option CYGIMP_POSIX_MQUEUE_VALIDATE_DESCRIPTOR {
            display          "Validate queue descriptors"
            flavor           bool
            default_value    1
            description      "
                This option turns on checking that message queue descriptors
                (of type mqd_t) passed into mq_* functions are valid. If so,
                the functions will fail with EBADF, as POSIX 1003.1 mandates.
                If this option is disabled, if an invalid descriptor is used,
                random corruption may occur, or the system may crash. If
                you are confident invalid descriptors will not be used,
                you may wish to be disable this to save some per-instance
                memory and execution time."
        }

        cdl_option CYGFUN_POSIX_MQUEUE_NOTIFY {
            display          "Allow empty queue notification"
            flavor           bool
            requires         CYGPKG_POSIX_SIGNALS
            default_value    CYGPKG_POSIX_SIGNALS
            description      "
                Enabling this option adds the function mq_notify() to the
                API. Without it, some code and per-message queue descriptor
                space is saved, as well as no longer requiring POSIX realtime
                signal support."
        }
    }

    # ----------------------------------------------------------------
    # Signals component

    cdl_component CYGPKG_POSIX_SIGNALS {
	display          "POSIX signals configuration"
	flavor           bool
	default_value    1
	requires	 CYGPKG_KERNEL_EXCEPTIONS
        requires         CYGPKG_POSIX_PTHREAD
        requires         CYGPKG_POSIX_TIMERS
        implements       CYGINT_POSIX_REALTIME_SIGNALS
        implements       CYGINT_ISO_SIGSETJMP
        requires         { CYGBLD_ISO_SIGSETJMP_HEADER == \
                             "<cyg/posix/sigsetjmp.h>" }
        implements       CYGINT_ISO_SIGNAL_NUMBERS
        implements       CYGINT_ISO_SIGNAL_IMPL
        requires         { CYGBLD_ISO_SIGNAL_NUMBERS_HEADER == \
                             "<cyg/posix/signal.h>" }
        requires         { CYGBLD_ISO_SIGNAL_IMPL_HEADER == \
                             "<cyg/posix/signal.h>" }
	description      "This component provides configuration controls for
	                  the POSIX signals."
        compile          signal.cxx except.cxx 
    }

    # ----------------------------------------------------------------
    # uname structure component

    cdl_component CYGPKG_POSIX_UTSNAME {
	display           "POSIX utsname configuration"
	flavor            bool
	default_value     1
	requires          { CYGBLD_ISO_UTSNAME_HEADER == \
                            "<cyg/posix/utsname.h>" }
	description       "This component provides configuration controls for
	                   the POSIX utsname structure and the uname() function."

	cdl_option CYG_POSIX_UTSNAME_LENGTH {
	    display          "Length of name strings in utsname structure"
	    flavor           data
	    default_value    65
	    legal_values     1 to 99999999
	}

	cdl_option CYG_POSIX_UTSNAME_NODENAME_LENGTH {
	    display          "Length of nodename string in utsname structure"
	    flavor           data
	    default_value    { CYG_POSIX_UTSNAME_LENGTH }
	    legal_values     1 to 99999999	    
	}

    }

    # ----------------------------------------------------------------
    # Tests

        cdl_option CYGPKG_POSIX_TESTS {
            display "POSIX tests"
            flavor  data
            no_define
            calculated { "tests/pthread1 tests/pthread2 tests/pthread3 tests/mutex3 tests/signal1 tests/timer1 tests/tm_basic tests/signal2 tests/mqueue1 tests/mqueue2 tests/sigsetjmp" }
            description   "
                This option specifies the set of tests for the POSIX package."
        }

}

# ====================================================================
# End of posix.cdl


