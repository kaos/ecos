# ====================================================================
##
##      hal_cortexm_ek_lm3s811.cdl
##
##      Stellaris Cortex-M3 EK-LM3S811 board platform HAL
##
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2011 Free Software Foundation, Inc.                        
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      ccoutand
# Contributors:   
# Date:           2011-01-18
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_CORTEXM_EK_LM3S811 {
    display       "Stellaris EK-LM3S811 Development Board HAL"
    doc           ref/hal-cortexm-lm3s-ek_lm3s811.html
    parent        CYGPKG_HAL_CORTEXM_LM3S8XX
    define_header hal_cortexm_ek_lm3s811.h
    include_dir   cyg/hal
    hardware

    description   "
        The EK-LM3S811 HAL package provides the support needed to run
        eCos on the Stellaris EK-LM3S811 EVAL board."

    compile       ek_lm3s811_misc.c platform_i2c.c

    requires      { CYGHWR_HAL_CORTEXM_LM3S == "LM3S8XX" }
    requires      { CYGHWR_HAL_CORTEXM_LM3S8XX == "LM3S811" }
    requires      { CYGNUM_HAL_CORTEXM_LM3S8XX_XTAL_FREQ == 6000000 }
    requires      { CYGHWR_HAL_CORTEXM_LM3S8XX_CLOCK_EXT == 1 }

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_cortexm_ek_lm3s811.h>"
        puts $::cdl_header "#include <pkgconf/hal_cortexm_lm3s8xx.h>"
        puts $::cdl_header "#define HAL_PLATFORM_CPU    \"Cortex-M3 - LM3S811\""
        puts $::cdl_header "#define HAL_PLATFORM_BOARD  \"Stellaris EK-LM3S811\""
        puts $::cdl_header "#define HAL_PLATFORM_EXTRA  \"\""
    }
}

# EOF hal_cortexm_ek_lm3s811.cdl
