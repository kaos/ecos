# ====================================================================
#
#      ser_arm_lpc24xx.cdl
#
#      eCos serial ARM/LPC24XX configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
## Copyright (C) 2004 eCosCentric Limited 
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Uwe Kindler  
# Original data:  gthomas, jskov
# Contributors:
# Date:           2008-07-06
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_IO_SERIAL_ARM_LPC24XX {
    display       "ARM LPC24xx serial device drivers"

    parent        CYGPKG_IO_SERIAL_DEVICES
    active_if     CYGPKG_IO_SERIAL
    active_if     CYGPKG_HAL_ARM_LPC24XX
    implements    CYGINT_IO_SERIAL_GENERIC_16X5X_CHAN_INTPRIO
    requires      CYGPKG_ERROR
    include_dir   cyg/io

    description   "
           This option enables the serial device drivers for the
           ARM LPC24xx."

    # FIXME: This really belongs in the GENERIC_16X5X package
    cdl_interface CYGINT_IO_SERIAL_GENERIC_16X5X_REQUIRED {
        display   "Generic 16x5x serial driver required"
    }
    define_proc {
        puts $::cdl_header "#define CYGPRI_IO_SERIAL_GENERIC_16X5X_STEP 4"
    }


    define_proc {
        puts $::cdl_system_header "/***** serial driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_GENERIC_16X5X_INL <cyg/io/arm_lpc24xx_ser.inl>"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_GENERIC_16X5X_CFG <pkgconf/io_serial_arm_lpc24xx.h>"
        puts $::cdl_system_header "/*****  serial driver proc output end  *****/"
    }
    
    # Support up to 4 on-chip UART modules. The number may vary between
    # processor variants so it is easy to update this here
    for { set ::channel 0 } { $::channel < 4 } { incr ::channel } {
    
        cdl_interface CYGINT_IO_SERIAL_LPC24XX_UART[set ::channel] {
            display     "Platform provides UART [set ::channel]"
            flavor      bool
            description "
                This interface will be implemented if the specific LPC24xx
                processor being used has on-chip UART [set ::channel], and if
                that UART is accessible on the target hardware."
        }

        cdl_component CYGPKG_IO_SERIAL_ARM_LPC24XX_SERIAL[set ::channel] {
            display       "ARM LPC24cxx UART [set ::channel] driver"
            flavor        bool
            active_if     CYGINT_IO_SERIAL_LPC24XX_UART[set ::channel]
            default_value 1

           implements CYGINT_IO_SERIAL_GENERIC_16X5X_REQUIRED
           implements CYGINT_IO_SERIAL_FLOW_CONTROL_HW
           implements CYGINT_IO_SERIAL_LINE_STATUS_HW

           description   "
                This option includes the serial device driver for the ARM
                LPC24xx UART [set ::channel]."

            cdl_option CYGDAT_IO_SERIAL_ARM_LPC24XX_SERIAL[set ::channel]_NAME {
                display       "Device name for UART [set ::channel]"
                flavor        data
                default_value   [format {"\"/dev/ser%d\""} $::channel]
                description   "
                    This option specifies the name of the serial device
                    for the ARM LPC24xx UART [set ::channel]."
            }

            cdl_option CYGNUM_IO_SERIAL_ARM_LPC24XX_SERIAL[set ::channel]_BAUD {
                display       "Baud rate for UART [set ::channel]"
                flavor        data
                legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 
                                2400 3600 4800 7200 9600 14400 19200 38400
                                57600 115200 230400 }
                default_value 38400
                description   "
                    This option specifies the default baud rate (speed)
                    for the ARM LPC24xx UART [set ::channel]."
            }

            cdl_option CYGNUM_IO_SERIAL_ARM_LPC24XX_SERIAL[set ::channel]_BUFSIZE {
                display       "Buffer size for the UART [set ::channel]"
                flavor        data
                legal_values  0 to 8192
                default_value 128
                description   "
                    This option specifies the size of the internal buffers
                    used for the ARM LPC24xx UART [set ::channel]."
            }
            
            cdl_option CYGNUM_IO_SERIAL_ARM_LPC24XX_SERIAL[set ::channel]_INTPRIO {
                display       "Interrupt priority of UART [set ::channel]"
                flavor        data
                legal_values  0 to 15
                default_value 15
                description   "
                    This option selects the interupt priority for the
                    UART [set ::channel] interrupts. There are 16
                    priority levels corresponding to the values 0
                    through 15 decimal, of which 15 is the lowest
                    priority. The reset value of these registers
                    defaults all interrupt to the lowest priority,
                    allowing a single write to elevate the priority of
                    an individual interrupt."
            }
        }
    }

     cdl_component CYGPKG_IO_SERIAL_ARM_LPC24XX_TESTING {
        display    "Testing parameters"
        flavor     bool
        calculated 1
        active_if  CYGPKG_IO_SERIAL_ARM_LPC24XX_SERIAL0

        implements CYGINT_IO_SERIAL_TEST_SKIP_9600
        implements CYGINT_IO_SERIAL_TEST_SKIP_115200
        implements CYGINT_IO_SERIAL_TEST_SKIP_PARITY_EVEN
        
        cdl_option CYGPRI_SER_TEST_SER_DEV {
            display       "Serial device used for testing"
            flavor        data
            default_value { CYGDAT_IO_SERIAL_ARM_LPC24XX_SERIAL0_NAME }
        }

        define_proc {
            puts $::cdl_header "#define CYGPRI_SER_TEST_CRASH_ID \"armlpc24xx\""
            puts $::cdl_header "#define CYGPRI_SER_TEST_TTY_DEV  \"/dev/tty0\""
        }
    }
}

# EOF ser_arm_lpc24xx.cdl
