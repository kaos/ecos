# ====================================================================
#
#      ser_i386_pc.cdl
#
#      eCos serial PC configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      nickg
# Original data:  gthomas, jskov, pjo
# Contributors:
# Date:           2000-02-14
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_component CYGPKG_IO_SERIAL_I386_PC_SERIAL0 {
    display       "PC serial port 0 driver"
    flavor        bool
    default_value 0
    description   "
        This option includes the serial device driver for port 0 on the 
        PC."

    cdl_option CYGDAT_IO_SERIAL_I386_PC_SERIAL0_NAME {
        display       "Device name for PC serial port 0"
        flavor        data
        default_value {"\"/dev/ser0\""}
        description   "
            This option specifies the device name port 0 on the PC."
    }

    cdl_option CYGNUM_IO_SERIAL_I386_PC_SERIAL0_BAUD {
        display       "Baud rate for the PC serial port 0 driver"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 234000
        }
        default_value 38400
        description   "
            This option specifies the default baud rate (speed) for the
            PC port 0."
    }

    cdl_option CYGNUM_IO_SERIAL_I386_PC_SERIAL0_BUFSIZE {
        display       "Buffer size for the PC serial port 0 driver"
        flavor        data
        legal_values  0 to 8192
        default_value 128
        description   "
            This option specifies the size of the internal buffers used
            for the PC port 0."
    }

    cdl_option CYGNUM_IO_SERIAL_I386_PC_SERIAL0_IOBASE {
	display "I/O base address for the i386-PC serial port 0"
	flavor    data
	legal_values 0 to 0xFF8
	default_value 0x3F8
	description "
	This option specifies the I/O address of the 8250 or 16550 for serial port 0."
    }

    cdl_option CYGNUM_IO_SERIAL_I386_PC_SERIAL0_IRQ {
	display "IRQ for the i386-PC serial port 0"
	flavor    data
	legal_values 0 to 15
	default_value 4
	description "
	This option specifies the IRQ of the 8250 or 16550 for serial port 0."
   }

    cdl_option CYGNUM_IO_SERIAL_I386_PC_SERIAL0_INT {
	display "IRQ for the i386-PC serial port 0"
	flavor    data
	legal_values 32 to 47
	default_value { CYGNUM_IO_SERIAL_I386_PC_SERIAL0_IRQ + 32 }
	description "
	This option specifies the interrupt vector of the 8250 or 16550 for serial port 0."
   }
}

cdl_component CYGPKG_IO_SERIAL_I386_PC_SERIAL1 {
    display       "PC serial port 1 driver"
    flavor        bool
    default_value 0
    description   "
        This option includes the serial device driver for port 1 on
        the PC."

    cdl_option CYGDAT_IO_SERIAL_I386_PC_SERIAL1_NAME {
        display       "Device name for PC serial port 1"
        flavor        data
        default_value {"\"/dev/ser1\""}
        description   "
            This option specifies the device name port 1 on the PC."
    }

    cdl_option CYGNUM_IO_SERIAL_I386_PC_SERIAL1_BAUD {
        display       "Baud rate for the PC serial port 1 driver"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 234000
        }
        default_value 38400
        description   "
            This option specifies the default baud rate (speed) for the
	    PC port 1."
    }

    cdl_option CYGNUM_IO_SERIAL_I386_PC_SERIAL1_BUFSIZE {
        display       "Buffer size for the PC serial port 1 driver"
        flavor        data
        legal_values  0 to 8192
        default_value 128
        description   "
            This option specifies the size of the internal buffers used
	    for the PC port 1."
    }

    cdl_option CYGNUM_IO_SERIAL_I386_PC_SERIAL1_IOBASE {
	display "I/O base address for the i386-PC serial port 1"
	flavor    data
	legal_values 0 to 0xFF8
	default_value 0x2F8
	description "
	This option specifies the I/O address of the 8250 or 16550 for serial port 1."
    }

    cdl_option CYGNUM_IO_SERIAL_I386_PC_SERIAL1_IRQ {
	display "IRQ for the i386-PC serial port 1"
	flavor    data
	legal_values 0 to 15
	default_value 3
	description "
	This option specifies the IRQ of the 8250 or 16550 for serial port 1."
   }

    cdl_option CYGNUM_IO_SERIAL_I386_PC_SERIAL1_INT {
	display "IRQ for the i386-PC serial port 1"
	flavor    data
	legal_values 32 to 47
	default_value { CYGNUM_IO_SERIAL_I386_PC_SERIAL1_IRQ + 32 }
	description "
	This option specifies the interrupt vector of the 8250 or 16550 for serial port 1."
   }
}
