# ====================================================================
#
#      io_pci.cdl
#
#      eCos PCI library configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Contributors:
# Date:           1999-08-12
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_IO_PCI {
    display       "PCI configuration library"
    doc           redirect/ecos-device-drivers.html
    include_dir   cyg/io
    parent        CYGPKG_IO
    description   "
           The PCI configuration library provides initialization of devices
           on the PCI bus. Functions to find and access these devices are
	   also provided."

    compile       pci.c pci_hw.c

    cdl_component CYGPKG_IO_PCI_OPTIONS {
        display "PCI build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_IO_PCI_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the PCI configuration library. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_IO_PCI_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the PCI configuration library. These flags are removed from
                the set of global flags if present."
        }

        cdl_option CYGPKG_IO_PCI_DEBUG {
            display "Enable debugging."
            flavor  bool
            default_value 0
            description   "
                This option enables minimal debugging of the PCI library.
                In particular, it will print information about devices as the
                PCI bus is being scanned/searched."
        }

        cdl_option CYGPKG_IO_PCI_TESTS {
            display "PCI tests"
            flavor  data
            no_define
            calculated { "tests/pci1 tests/pci2" }
            description   "
                This option specifies the set of tests for the PCI configuration library."
        }
    }
}
