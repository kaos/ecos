# ====================================================================
#
#      libc.cdl
#
#      C library configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      bartv
# Original data:  jlarmour
# Contributors:
# Date:           1999-06-13
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_LIBC {
    display       "C library"
    description   "
        This package enables compatibility with the ISO
        C standard - ISO/IEC 9899:1990. This allows the
        user application to use well known standard
        C library functions, and in eCos starts a
        thread to invoke the user function main()"
    doc           redirect/the-iso-standard-c-and-math-libraries.html
    compile       ctype/isalnum.cxx ctype/isalpha.cxx   ctype/iscntrl.cxx    \
                  ctype/isdigit.cxx ctype/isgraph.cxx   ctype/islower.cxx    \
                  ctype/isprint.cxx ctype/ispunct.cxx   ctype/isspace.cxx    \
                  ctype/isupper.cxx ctype/isxdigit.cxx  ctype/tolower.cxx    \
                  ctype/toupper.cxx                                          \
                                                                             \
                  errno/errno.cxx                                            \
                                                                             \
                  i18n/locale.cxx                                            \
                                                                             \
                  setjmp/longjmp.cxx                                         \
                                                                             \
                  signal/raise.cxx              signal/siginit.cxx           \
                  signal/signal.cxx                                          \
                                                                             \
                  stdio/common/fclose.cxx       stdio/common/fflush.cxx      \
                  stdio/common/fopen.cxx        stdio/common/freopen.cxx     \
                  stdio/common/setvbuf.cxx      stdio/common/snprintf.cxx    \
                  stdio/common/sprintf.cxx      stdio/common/sscanf.cxx      \
                  stdio/common/stderr.cxx       stdio/common/stdin.cxx       \
                  stdio/common/stdiofiles.cxx                                \
                  stdio/common/stdioinlines.cxx stdio/common/stdiosupp.cxx   \
                  stdio/common/stdout.cxx       stdio/common/stream.cxx      \
                  stdio/common/streambuf.cxx    stdio/common/ungetc.cxx      \
                  stdio/common/vsnprintf.cxx    stdio/common/vsscanf.cxx     \
                  stdio/input/fgetc.cxx         stdio/input/fgets.cxx        \
                  stdio/input/fread.cxx         stdio/input/fscanf.cxx       \
                  stdio/input/gets.cxx          stdio/input/scanf.cxx        \
                  stdio/input/vfscanf.cxx       stdio/output/fnprintf.cxx    \
                  stdio/output/fprintf.cxx      stdio/output/fputc.cxx       \
                  stdio/output/fputs.cxx        stdio/output/fwrite.cxx      \
                  stdio/output/printf.cxx       stdio/output/vfnprintf.cxx   \
                                                                             \
                  stdlib/_exit.cxx   stdlib/abort.cxx    stdlib/abs.cxx      \
                  stdlib/atexit.cxx  stdlib/atof.cxx     stdlib/atoi.cxx     \
                  stdlib/atol.cxx    stdlib/bsearch.cxx  stdlib/div.cxx      \
                  stdlib/exit.cxx    stdlib/getenv.cxx   stdlib/itoa.cxx     \
                  stdlib/labs.cxx    stdlib/ldiv.cxx     stdlib/malloc.cxx   \
                  stdlib/qsort.cxx   stdlib/rand.cxx     stdlib/strtod.cxx   \
                  stdlib/strtol.cxx  stdlib/strtoul.cxx  stdlib/system.cxx   \
                                                                             \
                  string/memchr.cxx  string/memcmp.cxx  string/memmove.cxx   \
                  string/strcat.cxx  string/strchr.cxx  string/strcmp.cxx    \
                  string/strcoll.cxx string/strcpy.cxx  string/strcspn.cxx   \
                  string/strlen.cxx  string/strncat.cxx string/strncmp.cxx   \
                  string/strncpy.cxx string/strpbrk.cxx string/strrchr.cxx   \
                  string/strspn.cxx  string/strstr.cxx  string/strsuppt.cxx  \
                  string/strtok.cxx  string/strxfrm.cxx                      \
                                                                             \
                  support/cstartup.cxx           support/environ.cxx         \
                  support/invokemain.cxx         support/main.cxx            \
                  support/mainthread.cxx                                     \
                                                                             \
                  time/asctime.cxx     time/asctime_r.cxx time/clock.cxx     \
                  time/ctime.cxx       time/ctime_r.cxx   time/difftime.cxx  \
                  time/gmtime.cxx      time/gmtime_r.cxx  time/localtime.cxx \
                  time/localtime_r.cxx time/mktime.cxx    time/settime.cxx   \
                  time/strftime.cxx    time/time.cxx      time/timeutil.cxx
    

    cdl_option CYGIMP_LIBC_CTYPE_INLINES {
        display       "Inline versions of <ctype.h> functions"
        default_value 1
        description   "
            This option chooses whether the simple character
            classification and conversion functions (e.g.
            isupper(), isalpha(), toupper(), etc.)
            from <ctype.h> are available as inline
            functions. This may improve performance and as
            the functions are small, may even improve code
            size."
    }

    # STRING CONFIGURATION OPTIONS
    cdl_component CYGPKG_LIBC_STRING {
        display       "String functions"
        flavor        none
        description   "
            Options associated with the standard string functions"

        script        string.cdl
    }

    # SETJMP CONFIGURATION OPTIONS
    cdl_option CYGIMP_LIBC_SETJMP_INLINES {
        display       "Inline version of the longjmp() function"
        default_value 1
        description   "
            This option chooses whether the longjmp() function
            is available as an inline function. This may
            improve performance, and as the function is small
            may even improve code size. "
    }

    # STDLIB CONFIGURATION OPTIONS
    cdl_component CYGPKG_LIBC_STDLIB {
        display       "Standard utility functions"
        flavor        none
        description   "
            Options associated with the standard utility functions in <stdlib.h>"

        script        stdlib.cdl
    }

    # STDIO CONFIGURATION OPTIONS
    cdl_component CYGPKG_LIBC_STDIO {
        display       "Standard input/output functions"
        flavor        bool
        requires      CYGPKG_IO
        requires      CYGPKG_IO_SERIAL_HALDIAG
        default_value 1
        description   "
            This enables support for standard I/O functions from <stdio.h>."

        script        stdio.cdl
    }


    # INTERNATIONALIZATION AND LOCALIZATION OPTIONS
    cdl_option CYGNUM_LIBC_MAX_LOCALE_NAME_SIZE {
        display       "Size of locale name strings"
        flavor        data
        legal_values  2 to 0x7fffffff
        default_value 16
        description   "
            This option controls the maximum size of
            locale names and is used, among other things
            to instantiate a static string used
            as a return value from the
            setlocale() function. When requesting the
            current locale settings with LC_ALL, a string
            must be constructed to contain this data, rather
            than just returning a constant string. This
            string data is stored in the static string.
            This depends on the length of locale names,
            hence this option. If just the C locale is
            present, this option can be set as low as 2."
    }

    # SIGNAL CONFIGURATION OPTIONS
    cdl_component CYGPKG_LIBC_SIGNALS {
        display       "Signals"
        flavor        bool
        default_value 1
        description   "
            This component controls signal functionality,
            as implemented in ISO C chapter 7.7 with the
            signal() and raise() functions. As well as
            allowing a program to send itself signals, it is
            also possible to cause hardware exceptions to
            be signalled to the program in a similar way."
        
        script        signals.cdl
    }


    # STARTUP OPTIONS
    cdl_component CYGPKG_LIBC_STARTUP {
        display       "ISO C startup/termination"
        flavor        none
        doc           redirect/c-library-startup.html
        description   "
            This component manages the control of the
            environment (in the general sense) that the
            C library provides for use for full ISO C
            compatibility, including a main() entry point
            supplied with arguments and an environment
            (as retrievable by the getenv() function).
            It also includes at the other end of things,
            what happens when main() returns or exit() is
            called."

        script        startup.cdl
    }

    # ERRNO OPTIONS
    cdl_component CYGPKG_LIBC_ERRNO {
        display       "errno"
        flavor        none
        description   "
            This package controls the behaviour of the
            errno variable (or more strictly, expression)
            from <errno.h>."

        cdl_option CYGSEM_LIBC_PER_THREAD_ERRNO {
            display       "Per-thread errno"
            requires      CYGVAR_KERNEL_THREADS_DATA
            default_value 1
            description   "
                This option controls whether the standard error
                code reporting variable errno is a per-thread
                variable, rather than global. Enabling this
                option will use one slot of kernel per-thread data.
                You should ensure you have enough slots configured
                for all your per-thread data."
        }

        cdl_option CYGNUM_LIBC_ERRNO_TRACE_LEVEL {
            display       "Tracing level"
            flavor        data
            legal_values  0 to 1
            default_value 0
            description   "
                Trace verbosity level for debugging the errno
                retrieval mechanism in errno.cxx. Increase this
                value to get additional trace output."
        }
    }

    # TIME OPTIONS
    cdl_component CYGPKG_LIBC_TIME {
        display       "Date/time"
        flavor        none
        description   "
            Options for date and time related functions from <time.h>"

        script        time.cdl
    }

    define_proc {
        puts $::cdl_header "/***** proc output start *****/"
        puts $::cdl_header "#include <pkgconf/system.h>"

        # MISCELLANEOUS DEFINES
        # These are not really adjustable by the user. Do not change these unless
        # you know what you are doing!

        # How to define inline functions
        puts $::cdl_header "#define CYGPRI_LIBC_INLINE extern __inline__"

        # The following isn't supported yet - I'm leaving it for now
        puts $::cdl_header "#ifdef __GNUC__xxxxxx"
        puts $::cdl_header "# define CYGPRI_LIBC_ATTRIB_FORMAT_STRFTIME __attribute__ ((format (strftime, 3)))"
        puts $::cdl_header "#else"
        puts $::cdl_header "# define CYGPRI_LIBC_ATTRIB_FORMAT_STRFTIME"
        puts $::cdl_header "#endif"

        # The following are only for compatibility, and will
        # eventually be removed once they are eliminated entirely from
        # the code base
        puts $::cdl_header "#define CYGPRI_LIBC_WEAK CYGBLD_ATTRIB_WEAK"

        # How to define aliases
        puts $::cdl_header "#define CYGPRI_LIBC_ALIAS(__symbol__) __attribute__ ((alias (__symbol__)))"

        puts $::cdl_header "# define CYGPRI_LIBC_WEAK_ALIAS(__symbol__) CYGBLD_ATTRIB_WEAK CYGPRI_LIBC_ALIAS(__symbol__)"

        # How to define functions that don't return
        puts $::cdl_header "#define CYGPRI_LIBC_NORETURN CYGBLD_ATTRIB_NORET"
        puts $::cdl_header "/****** proc output end ******/"
    }

    cdl_component CYGPKG_LIBC_OPTIONS {
        display "C library build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_LIBC_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the C library. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_LIBC_CFLAGS_REMOVE {
            display "Supressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the C library. These flags are removed from
                the set of global flags if present."
        }

        cdl_option CYGPKG_LIBC_TESTS {
            display "C library tests"
            flavor  data
            no_define
            calculated { "tests/ctype/ctype tests/i18n/setlocale tests/setjmp/setjmp tests/signal/signal1 tests/signal/signal2 tests/stdio/sprintf1 tests/stdio/sprintf2 tests/stdio/sscanf tests/stdio/stdiooutput tests/stdlib/abs tests/stdlib/atexit tests/stdlib/atoi tests/stdlib/atol tests/stdlib/bsearch tests/stdlib/div tests/stdlib/getenv tests/stdlib/labs tests/stdlib/ldiv tests/stdlib/qsort tests/stdlib/malloc1 tests/stdlib/malloc2 tests/stdlib/malloc3 tests/stdlib/rand1 tests/stdlib/rand2 tests/stdlib/rand3 tests/stdlib/rand4 tests/stdlib/realloc tests/stdlib/srand tests/stdlib/strtol tests/stdlib/strtoul tests/string/memchr tests/string/memcmp1 tests/string/memcmp2 tests/string/memcpy1 tests/string/memcpy2 tests/string/memmove1 tests/string/memmove2 tests/string/memset tests/string/strcat1 tests/string/strcat2 tests/string/strchr tests/string/strcmp1 tests/string/strcmp2 tests/string/strcoll1 tests/string/strcoll2 tests/string/strcpy1 tests/string/strcpy2 tests/string/strcspn tests/string/strcspn tests/string/strlen tests/string/strncat1 tests/string/strncat2 tests/string/strncpy1 tests/string/strncpy2 tests/string/strpbrk tests/string/strrchr tests/string/strspn tests/string/strstr tests/string/strtok tests/string/strxfrm1 tests/string/strxfrm2 tests/time/asctime tests/time/clock tests/time/ctime tests/time/gmtime tests/time/localtime tests/time/mktime tests/time/strftime tests/time/time" }
            description   "
                This option specifies the set of tests for the C library."
        }
    }
}
