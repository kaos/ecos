# ====================================================================
#
#      hal_sh_sh7750_dreamcast.cdl
#
#      SEGA Dreamcast HAL package configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      t@keshi.org
# Contributors:   t@keshi.org, jskov
# Date:           2001-07-30
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_SH_SH7750_DREAMCAST {
    display       "SEGA Dreamcast"
    parent        CYGPKG_HAL_SH
    requires      CYGPKG_HAL_SH_7750
    requires      ! CYGHWR_HAL_SH_BIGENDIAN
    define_header hal_sh_sh7750_dreamcast.h
    include_dir   cyg/hal
    description   "
        The HAL package provides the support needed to run
        eCos on SEGA Dreamcast."

    requires      { is_active(CYGSEM_REDBOOT_SH_LINUX_BOOT) implies 
                       (CYGDAT_REDBOOT_SH_LINUX_BOOT_ENTRY == 0x8c210000) }
    requires      { is_active(CYGSEM_REDBOOT_SH_LINUX_BOOT) implies 
                       (CYGDAT_REDBOOT_SH_LINUX_BOOT_BASE_ADDR == 0x8c001000) }
    requires      { is_active(CYGSEM_REDBOOT_SH_LINUX_BOOT) implies 
                       (CYGDAT_REDBOOT_SH_LINUX_BOOT_COMMAND_LINE == "mem=16M") }

    compile       hal_diag.c plf_misc.c dreamcast_pci.c fb_support.c
    compile       -library=libextras.a boot.S

    implements    CYGINT_HAL_DEBUG_GDB_STUBS
    implements    CYGINT_HAL_DEBUG_GDB_STUBS_BREAK
    implements    CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT
    implements    CYGINT_HAL_PLF_IF_INIT

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H   <pkgconf/hal_sh.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_sh_sh7750_dreamcast.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_IO_H <cyg/hal/plf_io.h>"
        puts $::cdl_header "#define CYGNUM_HAL_SH_SH4_SCIF_PORTS 1"
        puts $::cdl_header "#define CYGHWR_HAL_VSR_TABLE 0x8c010000"
        puts $::cdl_header "#define CYGHWR_HAL_VECTOR_TABLE 0x8c010100"
    }

    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        legal_values  {"RAM"}
        default_value {"RAM"}
        no_define
        define -file system.h CYG_HAL_STARTUP
        description   "
           When targetting the Dreamcast it is possible to build
           the system only for RAM bootstrap via a CD ROM."
    }

    cdl_option CYGSEM_DREAMCAST_FB_COMM {
        display        "Support framebuffer for communication channel"
        active_if      CYGPKG_REDBOOT
        flavor         bool
        default_value  1
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
        display      "Number of communication channels on the board"
        flavor       data
        calculated   1+CYGSEM_DREAMCAST_FB_COMM
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
        display          "Debug serial port"
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
           Dreamcast has only one serial port. This option
           chooses which port will be used to connect to a host
           running GDB."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
        display          "Diagnostic serial port"
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
           Dreamcast has only one serial port.  This option
           chooses which port will be used for diagnostic output."
    }

    cdl_option CYGNUM_HAL_SH_SH4_SCIF_BAUD_RATE_DEFAULT {
        flavor data
	calculated       115200
    };

    cdl_component CYGHWR_HAL_SH_PLF_CLOCK_SETTINGS {
        display          "SH on-chip platform clock controls"
        description      "
            The various clocks used by the system are derived from
            these options."
        flavor        none
        no_define
                     
        cdl_option CYGHWR_HAL_SH_OOC_XTAL {
            display          "SH clock crystal"
            flavor           data
            calculated       33333333
            no_define
            description      "
                This option specifies the frequency of the crystal all
                other clocks are derived from."
        }

        cdl_option CYGHWR_HAL_SH_OOC_CKIO {
            display          "SH clock CKIO output enable"
            default_value    1
            description      "
                This selects whether CKIO output is enabled."
        }

        cdl_option CYGHWR_HAL_SH_OOC_PLL_1 {
            display          "SH clock PLL circuit 1"
            flavor           data
            calculated       6
            description      "
                This selects whether PLL1 is enabled."
        }

        cdl_option CYGHWR_HAL_SH_OOC_PLL_2 {
            display          "SH clock PLL circuit 2"
            flavor           data
            calculated       1
            description      "
                This selects whether PLL2 is enabled."
        }

        cdl_option CYGHWR_HAL_SH_OOC_DIVIDER_1 {
            display          "SH clock first clock divider"
            flavor           data
            legal_values     { 1 2 }
            default_value    1
            no_define
            description      "
                First stage clock divider according to the mode (MD0..2).
                Set 2 for mode 2 and 4, otherwise set 1."
        }

        cdl_option CYGHWR_HAL_SH_OOC_DIVIDER_IFC {
            display          "SH clock divider, core"
            flavor           data
            calculated       1
            description      "
                This divider option affects the CPU core clock."
        }

        cdl_option CYGHWR_HAL_SH_OOC_DIVIDER_BFC {
            display          "SH clock divider, bus"
            flavor           data
            calculated       2
            description      "
                This divider option affects the bus clock."
        }

        cdl_option CYGHWR_HAL_SH_OOC_DIVIDER_PFC {
            display          "SH clock divider, peripheral"
            flavor           data
            calculated       4
            description      "
                This divider option affects the peripheral clock."
        }

        cdl_option CYGHWR_HAL_SH_OOC_CLOCK_MODE {
            display          "SH clock mode"
            flavor           data
            calculated       5
            description      "
                This option must mirror the clock mode hardwired on
                the MD0-MD2 pins of the CPU in order to correctly
                initialize the FRQCR register."
        }
    }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        parent  CYGPKG_NONE
        description   "
	    Global build options including control over
	    compiler flags, linker flags and choice of toolchain."


        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "sh-elf" }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { "-ml -m3 -Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -ggdb -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority" }
            description   "
                This option controls the global compiler flags which
                are used to compile all packages by
                default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { "-ml -m3 -ggdb -nostdlib -Wl,--gc-sections -Wl,-static" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }

        cdl_option CYGBLD_BUILD_GDB_STUBS {
            display "Build GDB stub ROM image"
            default_value 0
            requires CYGSEM_HAL_ROM_MONITOR
            requires CYGBLD_BUILD_COMMON_GDB_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT
            requires CYGDBG_HAL_DEBUG_GDB_THREAD_SUPPORT
            requires ! CYGDBG_HAL_COMMON_INTERRUPTS_SAVE_MINIMUM_CONTEXT
            requires ! CYGDBG_HAL_COMMON_CONTEXT_SAVE_MINIMUM
            no_define
            description "
                This option enables the building of the GDB stubs for the
                board. The common HAL controls takes care of most of the
                build process, but the final conversion from ELF image to
                binary data is handled by the platform CDL, allowing
                relocation of the data if necessary."

            make -priority 320 {
                <PREFIX>/bin/gdb_module.bin : <PREFIX>/bin/gdb_module.img
                $(OBJCOPY) -O binary $< $@
            }
        }
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { "sh_sh7750_dreamcast_ram" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { "<pkgconf/mlt_sh_sh7750_dreamcast_ram.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { "<pkgconf/mlt_sh_sh7750_dreamcast_ram.h>" }
        }
    }

    cdl_option CYGSEM_HAL_USE_ROM_MONITOR {
        display       "Work with a ROM monitor"
        flavor        booldata
        legal_values  { "GDB_stubs" }
        default_value 0
        requires      { CYG_HAL_STARTUP == "RAM" }
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      !CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
        description   "
            Support can be enabled for boot ROMs or ROM monitors which contain
            GDB stubs. This support changes various eCos semantics such as
            the encoding of diagnostic output, and the overriding of hardware
            interrupt vectors."
    }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "ROM" }
        description   "
            Enable this option if this program is to be used as a ROM monitor,
            i.e. applications will be loaded into RAM on the board, and this
            ROM monitor may process exceptions or interrupts generated from the
            application. This enables features such as utilizing a separate
            interrupt stack when exceptions are generated."
    }
}
