# ====================================================================
#
#	iq80310_eth_drivers.cdl
#
#	Ethernet drivers
#	Intel IQ80310 and PRO/100+ platform specific support
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      hmt
# Original data:  hmt
# Contributors:	  gthomas
# Date:           2000-02-01
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_ARM_IQ80310 {
    display       "Intel IQ80310 with PRO/100+ ethernet driver"

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if     CYGPKG_IO_ETH_DRIVERS
    active_if     CYGPKG_HAL_ARM_IQ80310

    include_dir   cyg/io

    # FIXME: This really belongs in the INTEL_I82559 package
    cdl_interface CYGINT_DEVS_ETH_INTEL_I82559_REQUIRED {
        display   "Intel i82559 ethernet driver required"
    }

    define_proc {
        puts $::cdl_system_header "/***** ethernet driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_DEVS_ETH_INTEL_I82559_INL <cyg/io/devs_eth_iq80310.inl>"
        puts $::cdl_system_header "#define CYGDAT_DEVS_ETH_INTEL_I82559_CFG <pkgconf/devs_eth_arm_iq80310.h>"
        puts $::cdl_system_header "/*****  ethernet driver proc output end  *****/"
    }


    cdl_component CYGPKG_DEVS_ETH_ARM_IQ80310_ETH0 {
        display       "IQ80310 builtin ethernet port driver"
        flavor        bool
        default_value 1
        description   "
            This option includes the ethernet device driver for the
            IQ80310 builtin port."

        implements CYGHWR_NET_DRIVERS
        implements CYGHWR_NET_DRIVER_ETH0
        implements CYGINT_DEVS_ETH_INTEL_I82559_REQUIRED

        cdl_option CYGDAT_DEVS_ETH_ARM_IQ80310_ETH0_NAME {
            display       "Device name for the ETH0 ethernet port driver"
            flavor        data
            default_value {"\"eth0\""}
            description   "
                This option sets the name of the ethernet device for the
                IQ80310 builtin port."
        }

        cdl_option CYGNUM_DEVS_ETH_ARM_IQ80310_MAX_RX_DESCRIPTORS {
            display       "Maximum number of RX descriptors"
            flavor  data
            default_value { CYGPKG_REDBOOT ? 4 : 128 }
            define        MAX_RX_DESCRIPTORS
            description   "
                    An RX descriptor is used for each ethernet frame required
                    to be passed to the upper networking layers. This option
                    sets the maximum number of these. Higher numbers use more
                    memory, lower numbers will reduce performance. The system
                    appears to work OK with as few as 8 descriptors but limps
                    painfully with only 4. Performance is better with more than
                    8, but since the size of non-cached (so useless for anything
                    else) memory window is 1Mb, we might as well use it all.
                    128 RX and TX descriptors uses the whole 1Mb, near enough."
        }
    
        cdl_option CYGNUM_DEVS_ETH_ARM_IQ80310_MAX_TX_DESCRIPTORS {
            display       "Maximum number of TX descriptors"
            flavor  data
            default_value { CYGPKG_REDBOOT ? 4 : 128 }
            define        MAX_TX_DESCRIPTORS
            description   "
                    A TX descriptor is used for each ethernet frame passed down
                    from upper networking layers for transmission. This option
                    sets the maximum number of these. Higher numbers use more
                    memory, lower numbers will reduce performance. The system
                    appears to work OK with as few as 8 descriptors but limps
                    painfully with only 4. Performance is better with more than
                    8, but since the size of non-cached (so useless for anything
                    else) memory window is 1Mb, we might as well use it all.
                    128 RX and TX descriptors uses the whole 1Mb, near enough."
        }

        cdl_component CYGSEM_DEVS_ETH_ARM_IQ80310_ETH0_SET_ESA {
            display       "Set the ethernet station address"
            flavor        bool
	    default_value 0
            description   "Enabling this option will allow the ethernet
            station address to be forced to the value set by the
            configuration.  This may be required if the hardware does
            not include a serial EEPROM for the ESA."
            
            cdl_option CYGDAT_DEVS_ETH_ARM_IQ80310_ETH0_ESA {
                display       "The ethernet station address"
                flavor        data
                default_value {"{0x00, 0xB5, 0xE0, 0xB5, 0xE0, 0x11}"}
                description   "The ethernet station address"
            }
        }

    }

}

# EOF iq80310_eth_drivers.cdl
