# ====================================================================
#
#      i18n.cdl
#
#      C library internationalization (i18n) related configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jlarmour
# Contributors:
# Date:           2000-04-14
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_LIBC_I18N {
    display       "ISO C library internationalization functions"
    description   "
        This package provides internationalization functions specified by the
        ISO C standard - ISO/IEC 9899:1990. These include locale-related
        functionality and <ctype.h> functionality."
    doc           redirect/the-iso-standard-c-and-math-libraries.html
    include_dir   cyg/libc/i18n
    parent        CYGPKG_LIBC
    implements    CYGINT_ISO_LOCALE
    implements    CYGINT_ISO_CTYPE
    requires      CYGPKG_ISOINFRA
    compile       ctype.cxx locale.cxx

# ====================================================================

    cdl_option CYGNUM_LIBC_I18N_MAX_LOCALE_NAME_SIZE {
        display       "Size of locale name strings"
        flavor        data
        legal_values  2 to 0x7fffffff
        default_value 2
        description   "
            This option controls the maximum size of
            locale names and is used, among other things
            to instantiate a static string used
            as a return value from the
            setlocale() function. When requesting the
            current locale settings with LC_ALL, a string
            must be constructed to contain this data, rather
            than just returning a constant string. This
            string data is stored in the static string.
            This depends on the length of locale names,
            hence this option. If just the C locale is
            present, this option can be set as low as 2."
    }


# ====================================================================

    cdl_option CYGIMP_LIBC_I18N_CTYPE_INLINES {
        display       "Inline versions of <ctype.h> functions"
        default_value 1
        requires      { CYGBLD_ISO_CTYPE_HEADER == \
                           "<cyg/libc/i18n/ctype.inl>" }
        description   "
            This option chooses whether the simple character
            classification and conversion functions (e.g.
            isupper(), isalpha(), toupper(), etc.)
            from <ctype.h> are available as inline
            functions. This may improve performance and as
            the functions are small, may even improve code
            size."
    }

# ====================================================================

    cdl_component CYGPKG_LIBC_I18N_OPTIONS {
        display "C library i18n functions build options"
        flavor  none
        no_define
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_LIBC_I18N_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the C library. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_LIBC_I18N_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the C library. These flags are removed from
                the set of global flags if present."
        }

        cdl_option CYGPKG_LIBC_I18N_TESTS {
            display "C library i18n function tests"
            flavor  data
            no_define
            calculated { "tests/ctype tests/setlocale" }
            description   "
                This option specifies the set of tests for the C library
                i18n functions."
        }
    }
}

# ====================================================================
# EOF i18n.cdl
