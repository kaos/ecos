# ====================================================================
#
#      startup.cdl
#
#      C library startup related configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  jlarmour
# Contributors:
# Date:           1999-07-06
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_option CYGDAT_LIBC_ARGUMENTS {
    display       "Arguments to main()"
    flavor        data
    default_value {"{\"\", NULL}"}
    description   "
        This option allows the setting of the arguments
        to the main function. This only has any effect
        when cyg_iso_c_start() is used to start the
        ISO C compatibility. This will automatically
        invoke main() in an ISO C compatible fashion.
        This option is in fact used as argv, and so is
        an n-tuple of string constants. The final
        entry must be NULL. Conventionally if argv\[0\]
        is supplied, it is used to inform the program
        of its name."
}

cdl_component CYGSEM_LIBC_STARTUP_MAIN_THREAD {
    display       "main() invoked as thread"
    requires      CYGPKG_KERNEL
    flavor        bool
    default_value 1
    description   "
        It is normally expected (e.g. in a POSIX 1003.1
        environment) that main() is run in the context
        of a thread just like any other thread. If this
        option is disabled then main() will instead be
        called in the context of the initialization
        routines, without the scheduler running and
        using the interrupt stack. This means that 
        any functions that may require interactions
        with a running kernel will not work (including
        libc functions, if configured to be thread safe
        for example), so you should restrict yourself
        to only calling fully re-entrant functions from
        within main() in this case."

    cdl_component CYGSEM_LIBC_MAIN_STACK_FROM_SYSTEM {
        display        "System provides stack for main()'s thread"
        description    "
            This option controls whether the stack of
            main()'s thread is provided by the application or
            provided by the system. When disabled, the
            application must declare a pointer variable
            cyg_libc_main_stack which is a pointer to an
            appropriately aligned region of memory. The
            application must also declare a variable of
            type `int' called cyg_libc_main_stack_size
            which contains the size of the stack in bytes.
            This must be a multiple of 8."
        flavor         bool
        default_value  1

        cdl_option CYGNUM_LIBC_MAIN_DEFAULT_STACK_SIZE {
            display        "main()'s default thread stack size"
            flavor         data
            legal_values   16 to 0x7fffffff
            default_value  8192
            description    "
                With an eCos kernel, when the cyg_iso_c_start()
                function is used to invoke the user-supplied
                main() function in an ISO C compatible fashion,
                a separate thread is created to call main().
                This option controls the size of that thread's
                stack, which is allocated in the BSS. It
                must be a multiple of 8. Note, a low number
                here may be overriden by the HAL if there is
                a minimum requirement to process interrupts
                etc."
        }
    }

    cdl_option CYGNUM_LIBC_MAIN_THREAD_PRIORITY {
        display         "Priority of main()'s thread"
        description     "
            This option is used to provide the thread
            priority which main()'s thread runs at. Be
            sure to check that this number is appropriate
            for the kernel scheduler chosen. Different
            kernel schedulers impose different restrictions
            on the usable priorities."
        flavor          data
        legal_values    0 to 0x7fffffff
        default_value   10
   }
}

cdl_component CYGFUN_LIBC_ATEXIT {
    display        "Include atexit() function"
    flavor         bool
    default_value  1
    description    "
        This option enables the use of the atexit()
        function, and ensure that the atexit handlers
        are invoked from within exit() as defined in
        the ISO C standard."

    cdl_option CYGNUM_LIBC_ATEXIT_HANDLERS {
        display        "Number of functions atexit() supports"
        flavor         data
        legal_values   1 to 0x7fffffff
        default_value  32
        description    "
            This option sets the number of functions
            that atexit() has room for. In other words,
            the number of separate atexit() calls that
            can be made before calling exit() or returning
            from main() ( in an environment controlled by
            cyg_iso_c_start() ). For strict compliance
            with the ISO C standard this should be at
            least 32."
    }
}

cdl_option CYGSEM_LIBC_EXIT_CALLS_FFLUSH {
    display        "Make exit() call fflush()"
    requires       CYGSEM_LIBC_STDIO_WANT_BUFFERED_IO
    default_value  1
    description    "
        This option will ensure that all output
        streams are flushed when exitting using
        exit() as prescribed by the ISO C standard."
}

cdl_option CYGSEM_LIBC_EXIT_STOPS_SYSTEM {
    display        "_exit() stops all threads"
    requires       CYGPKG_KERNEL
    default_value  0
    description    "
        If this option is enabled then _exit(),
        which is called from exit() which itself is
        called on return from main(), stops the eCos
        scheduler. For strict POSIX 1003.1
        compatibility this would be the normal
        behaviour. To allow the thread to simply
        exit, without affecting other threads, simply
        disable this option. If there is no eCos
        scheduler, then _exit() simply loops
        irrespective of the setting of this option."
}

cdl_component CYGPKG_LIBC_ENVIRONMENT {
    display       "Provide a system environment"
    flavor         bool
    default_value  1
    description   "
        This option allows use of the getenv() function
        and the global environment pointer
        char **environ defined by POSIX 1003.1.
        Disabling this saves a small amount of space."

    cdl_option CYGDAT_LIBC_DEFAULT_ENVIRONMENT {
        display       "Default environment"
        flavor        data
        default_value {"{ NULL }"}
        description   "
            This option allows the setting of the default
            contents of the environment. This is in fact
            the contents of the global environment pointer
            char **environ defined by POSIX 1003.1. Strings
            must be of the form NAME=VALUE, and the final
            entry must be NULL."
    }
}

cdl_option CYGSEM_LIBC_INVOKE_DEFAULT_STATIC_CONSTRUCTORS {
    display        "Invoke default static constructors"
    requires       CYGSEM_HAL_STOP_CONSTRUCTORS_ON_FLAG
    requires       CYGSEM_LIBC_STARTUP_MAIN_THREAD
    default_value  0
    description    "
        This option causes the C library to call
        static constructors with default priority
        from within the context of the main() thread,
        working with the co-operation of the HAL.
        This may be needed for environments that
        expect static constructors to be run in a
        thread context. Note that this uses an object
        with priority 65534. Therefore do not use
        priority 65534 for any other static objects
        with this option enabled."
}
