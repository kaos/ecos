# ====================================================================
#
#      flash_bootblock.cdl
#
#      FLASH memory - Hardware support for Intel Boot Block Flash Memory
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
# -------------------------------------------
# This file is part of eCos, the Embedded Configurable Operating System.
# Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
#
# eCos is free software; you can redistribute it and/or modify it under
# the terms of the GNU General Public License as published by the Free
# Software Foundation; either version 2 or (at your option) any later version.
#
# eCos is distributed in the hope that it will be useful, but WITHOUT ANY
# WARRANTY; without even the implied warranty of MERCHANTABILITY or
# FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
# for more details.
#
# You should have received a copy of the GNU General Public License along
# with eCos; if not, write to the Free Software Foundation, Inc.,
# 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
#
# As a special exception, if other files instantiate templates or use macros
# or inline functions from this file, or you compile this file and link it
# with other works to produce a work based on this file, this file does not
# by itself cause the resulting work to be covered by the GNU General Public
# License. However the source code for this file must still be made available
# in accordance with section (3) of the GNU General Public License.
#
# This exception does not invalidate any other reasons why a work based on
# this file might be covered by the GNU General Public License.
#
# Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
# at http://sources.redhat.com/ecos/ecos-license
# -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Contributors:   jskov
# Date:           2000-07-26
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_FLASH_INTEL_BOOTBLOCK {
    display       "Intel boot block flash memory support"

    parent        CYGPKG_IO_FLASH
    active_if	  CYGPKG_IO_FLASH

    implements    CYGHWR_IO_FLASH_DEVICE
    implements    CYGHWR_IO_FLASH_DEVICE_NOT_IN_RAM

    include_dir   .
    include_files ; # none _exported_ whatsoever
    description   "FLASH memory device support for Intel boot block flash memory"
    compile       bootblock_flash.c

    make -priority 1 {
        flash_erase_block.o: $(REPOSITORY)/$(PACKAGE)/src/flash_erase_block.c
        $(CC) -S $(INCLUDE_PATH) $(CFLAGS) -g0 -mcpu=strongarm -fno-function-sections $(REPOSITORY)/$(PACKAGE)/src/flash_erase_block.c
        echo "#include <cyg/hal/arch.inc>" > flash_erase_block2.S
        cat  flash_erase_block.s >> flash_erase_block2.S
        echo "FUNC_END(flash_erase_block_end)" >>flash_erase_block2.S
        $(CC) -c $(INCLUDE_PATH) -o flash_erase_block.o flash_erase_block2.S
        $(AR) rcs $(PREFIX)/lib/libtarget.a flash_erase_block.o
    }
    make -priority 1 {
        flash_program_buf.o: $(REPOSITORY)/$(PACKAGE)/src/flash_program_buf.c
        $(CC) -S $(INCLUDE_PATH) $(CFLAGS) -g0 -mcpu=strongarm -fno-function-sections $(REPOSITORY)/$(PACKAGE)/src/flash_program_buf.c
        echo "#include <cyg/hal/arch.inc>" > flash_program_buf2.S
        cat  flash_program_buf.s >> flash_program_buf2.S
        echo "FUNC_END(flash_program_buf_end)" >>flash_program_buf2.S
        $(CC) -c $(INCLUDE_PATH) -o flash_program_buf.o flash_program_buf2.S
        $(AR) rcs $(PREFIX)/lib/libtarget.a flash_program_buf.o
    }
    make -priority 1 {
        flash_query.o: $(REPOSITORY)/$(PACKAGE)/src/flash_query.c
        $(CC) -S $(INCLUDE_PATH) $(CFLAGS) -g0 -mcpu=strongarm -fno-function-sections $(REPOSITORY)/$(PACKAGE)/src/flash_query.c
        echo "#include <cyg/hal/arch.inc>" > flash_query2.S
        cat  flash_query.s >> flash_query2.S
        echo "FUNC_END(flash_query_end)" >>flash_query2.S
        $(CC) -c $(INCLUDE_PATH) -o flash_query.o flash_query2.S
        $(AR) rcs $(PREFIX)/lib/libtarget.a flash_query.o
    }
}
