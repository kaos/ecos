# ====================================================================
#
#      flash_mips_qed_ocelot.cdl
#
#      FLASH memory - Hardware support for QED Ocelot board
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Contributors:   jskov
# Date:           2000-12-05
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_FLASH_MIPS_QED_OCELOT {
    display       "Flash memory support for QED Ocelot board"

    parent        CYGPKG_IO_FLASH
    active_if	  CYGPKG_IO_FLASH

    # FIXME: This really belongs in the ADM_AM29F040B package
    cdl_interface CYGINT_DEVS_FLASH_AMD_AM29F040B_REQUIRED {
        display   "AMD AM29F040B driver required"
    }

    include_dir   cyg/io
    description   "FLASH memory device support for QED Ocelot board"

    implements    CYGINT_DEVS_FLASH_AMD_AM29F040B_REQUIRED

    define_proc {
        puts $::cdl_system_header "/***** flash driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_DEVS_FLASH_AMD_AM29F040B_INL <cyg/io/devs_flash_mips_qed_ocelot.inl>"
        puts $::cdl_system_header "#define CYGDAT_DEVS_FLASH_AMD_AM29F040B_CFG <pkgconf/devs_flash_mips_qed_ocelot.h>"
        puts $::cdl_system_header "/*****  flash driver proc output end  *****/"
    }
}
