# ====================================================================
#
#      fatfs.cdl
#
#      FAT Filesystem configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 2003 Savin Zlobec 
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      savin 
# Contributors:   
# Date:           2003-06-25
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_FS_FAT {
    display         "FAT filesystem"
    include_dir     cyg/fatfs

    requires        CYGPKG_IO_FILEIO

    requires        CYGPKG_ISOINFRA
    requires        CYGINT_ISO_ERRNO
    requires        CYGINT_ISO_ERRNO_CODES
    requires        CYGPKG_MEMALLOC
    requires        CYGPKG_BLOCK_LIB
#    requires        CYGFUN_LIBC_STRING_BSD_FUNCS

    implements      CYGINT_IO_FILEIO_FS
    
    compile         -library=libextras.a fatfs.c        \
                                         fatfs_supp.c   \
                                         fatfs_ncache.c \
                                         fatfs_tcache.c

    cdl_option      CYGNUM_FS_FAT_NODE_HASH_TABLE_SIZE {
        display         "Node hash table size"
        flavor          data
        default_value   32
        legal_values    1 to 9999999999
        description     "This option controls the number of slots in the 
                         hash table used to store file nodes using filenames 
                         as keys."
    }

    cdl_option      CYGNUM_FS_FAT_NODE_ALLOC_THRESHOLD {
        display         "Node allocation treshold"
        flavor          data
        default_value   16
        legal_values    1 to 9999999999
        description     "This option controls at which point the filesystem 
                         starts reusing dead file nodes rather then allocating
                         memory for new nodes."
    }
   
    cdl_option      CYGNUM_FS_FAT_FAT_TABLE_CACHE_MEMSIZE {
        display         "FAT table cache memory size"
        flavor          data
        default_value   10240
        legal_values    1 to 9999999999
        description     "This option controls the amount of memory used
                         for the FAT table cache."
    }

    cdl_option      CYGNUM_FS_FAT_FAT_TABLE_CACHE_INCREMENT {
        display         "FAT table cache size increment"
        flavor          data
        default_value   10
        legal_values    1 to 9999999999
        description     "This option controls the amount of memory by which 
                         the per-file FAT table cache will grow."
    }
   
    cdl_option      CYGNUM_FS_FAT_BLOCK_CACHE_MEMSIZE {
        display         "FAT block cache memory size"
        flavor          data
        default_value   10240 
        legal_values    1 to 9999999999
        description     "This option controls the amount of memory used for 
                         the block cache."
    }

    cdl_option      CYGDBG_FS_FAT_NODE_CACHE_EXTRA_CHECKS {
        display         "Node cache extra checks"
        flavor          bool
        default_value   1
        active_if       CYGPKG_INFRA_DEBUG && CYGDBG_USE_ASSERTS
        description     "This option controls the inclusion of extra
                         sanity checks in node cache code."
    }
    
    # --------------------------------------------------------------------
    
    cdl_option      CYGPKG_FS_FAT_TESTS {
        display         "FAT FS tests"
        flavor          data
        no_define
        calculated      { "tests/fileio1.c" }
        description     "This option specifies the set of tests for the 
                         FAT FS package."
    }
}

# ====================================================================
# End of fatfs.cdl
