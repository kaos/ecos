# ====================================================================
#
#      romfs.cdl
#
#      ROM Filesystem configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2004, 2009 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      nickg
# Original data:  nickg
# Contributors:   richard.panton@3glab.com
# Date:           2000-08-01
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_FS_ROM {
    display        "ROM filesystem"
    doc            ref/fileio.html
    include_dir    cyg/romfs

    parent         CYGPKG_IO_FILEIO
    requires       CYGPKG_IO_FILEIO

    requires       CYGPKG_ISOINFRA
    requires       CYGINT_ISO_ERRNO
    requires       CYGINT_ISO_ERRNO_CODES

    implements     CYGINT_IO_FILEIO_FS
    
    compile        -library=libextras.a romfs.c

    cdl_option CYGBLD_FS_ROMFS_MK_ROMFS {
        display       "Build the tool used to build filesystems"
        flavor        bool
        default_value 1

        make -priority 98 {
            <PREFIX>/bin/file2c.tcl: <PACKAGE>/support/file2c.tcl
            @mkdir -p "$(dir $@)"
            @cp $< $@
        }

        # FIXME: host compiler/flags should be provided by config system
        make -priority 98 {
            <PREFIX>/bin/mk_romfs: <PACKAGE>/support/mk_romfs.c
            @mkdir -p "$(dir $@)"
            @$(HOST_CC) -g -O2 -o $@ $< || cc -g -O2 -o $@ $< || gcc -g -O2 -o $@ $<
        }

        description "
            When enabled this option will build a host tool which can be
            used to create a rom filesystem image."
    }

    cdl_option CYGPKG_FS_ROM_RET_DIRENT_DTYPE {
        display       "Support for fileio's struct dirent d_type field"
        flavor        bool
        default_value 0
        active_if     CYGPKG_FILEIO_DIRENT_DTYPE

        description "
            This option controls whether the ROM filesystem supports
            setting fileio's struct dirent d_type field.
            If this option is enabled, d_type will be set. Otherwise,
            nothing will be done, d_type's value will be zero because
            fileio already sets it."
    }

    # ----------------------------------------------------------------
    # Tests

    cdl_component CYGTST_ROMFS_BUILD_TESTS {
        display       "Build ROM filesystem tests"
        flavor        bool
        no_define
        default_value 0
        requires      CYGINT_LIBC_STARTUP_CONTEXT
        requires      CYGINT_ISO_STDIO_FORMATTED_IO
        requires      CYGINT_ISO_STRERROR
        requires      CYGBLD_FS_ROMFS_MK_ROMFS        
        description   "
                This option enables the building of the ROM filesystem tests."

        make -priority 100 {
            <PREFIX>/include/cyg/romfs/testromfs_le.h : <PACKAGE>/tests/testromfs <PREFIX>/bin/mk_romfs <PREFIX>/bin/file2c.tcl
            $(PREFIX)/bin/mk_romfs $< testromfs_le.bin
            @mkdir -p "$(dir $@)"
            tclsh $(PREFIX)/bin/file2c.tcl testromfs_le.bin $@
        }
    
        make -priority 100 {
            <PREFIX>/include/cyg/romfs/testromfs_be.h : <PACKAGE>/tests/testromfs <PREFIX>/bin/mk_romfs <PREFIX>/bin/file2c.tcl
            $(PREFIX)/bin/mk_romfs -b $< testromfs_be.bin
            @mkdir -p "$(dir $@)"
            tclsh $(PREFIX)/bin/file2c.tcl testromfs_be.bin $@
        }
    
        cdl_option CYGPKG_FS_ROM_TESTS {
            display "ROM filesystem tests"
            flavor  data
            no_define
            calculated { "tests/romfs1" }
                description   "
                    This option specifies the set of tests for the ROM filesystem package."
        }
    }
}

# End of romfs.cdl
