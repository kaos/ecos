# ====================================================================
#
#      ser_arm_cma230.cdl
#
#      eCos serial ARM/CMA230 configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  gthomas
# Contributors:
# Date:           1999-07-08
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_component CYGPKG_IO_SERIAL_ARM_CMA230_SERIAL_A {
    display       "Cogent ARM/CMA230 serial port A driver"
    flavor        bool
    default_value 0
    description   "
        This option includes the serial device driver for the Cogent 
        ARM/CMA230 port A."

    cdl_option CYGDAT_IO_SERIAL_ARM_CMA230_SERIAL_A_NAME {
        display       "Device name for Cogent ARM/CMA230 serial port A"
        flavor        data
        default_value {"\"/dev/ser1\""}
        description   "
            This option specifies the device name for the Cogent 
            ARM/CMA230 port A."
    }

    cdl_option CYGNUM_IO_SERIAL_ARM_CMA230_SERIAL_A_BAUD {
        display       "Baud rate for the Cogent ARM/CMA230 serial port A driver"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 234000
        }
        default_value 38400
        description   "
            This option specifies the default baud rate (speed) for the
            Cogent ARM/CMA230 port A."
    }

    cdl_option CYGNUM_IO_SERIAL_ARM_CMA230_SERIAL_A_BUFSIZE {
        display       "Buffer size for the Cogent ARM/CMA230 serial port A driver"
        flavor        data
        legal_values  0 to 8192
        default_value 128
        description   "
            This option specifies the size of the internal buffers used 
            for the Cogent ARM/CMA230 port A."
    }
}

cdl_component CYGPKG_IO_SERIAL_ARM_CMA230_SERIAL_B {
    display       "Cogent ARM/CMA230 serial port B driver"
    flavor        data
    default_value 0
    description   "
        This option includes the serial device driver for the Cogent 
        ARM/CMA230 port B."

    cdl_option CYGDAT_IO_SERIAL_ARM_CMA230_SERIAL_B_NAME {
        display       "Device name for Cogent ARM/CMA230 serial port B"
        flavor        data
        default_value {"\"/dev/ser2\""}
        description   "
            This option specifies the device name for the Cogent 
            ARM/CMA230 port B."
    }

    cdl_option CYGNUM_IO_SERIAL_ARM_CMA230_SERIAL_B_BAUD {
        display       "Baud rate for the Cogent ARM/CMA230 serial port B driver"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 234000
        }
        default_value 38400
        description   "
            This option specifies the default baud rate (speed) for the 
            Cogent ARM/CMA230 port B."
    }

    cdl_option CYGNUM_IO_SERIAL_ARM_CMA230_SERIAL_B_BUFSIZE {
        display       "Buffer size for the Cogent ARM/CMA230 serial port B driver"
        flavor        data
        legal_values  0 to 8192
        default_value 128
        description   "
            This option specifies the size of the internal buffers used 
            for the Cogent ARM/CMA230 port B."
    }
}
