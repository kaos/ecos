# ====================================================================
#
#      string.cdl
#
#      C library string related configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  jlarmour
# Contributors:
# Date:           1999-07-06
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_option CYGIMP_LIBC_STRING_INLINES {
    display       "Inline versions of <string.h> functions"
    default_value 1
    description   "
        This option chooses whether some of the
        particularly simple string functions from
        <string.h> are available as inline
        functions. This may improve performance, and as
        the functions are small, may even improve code
        size."
}

cdl_option CYGIMP_LIBC_STRING_PREFER_SMALL_TO_FAST {
    display       "Optimize string functions for code size"
    flavor bool
    default_value 0
    description   "
        This option tries to reduce string function
        code size at the expense of execution speed. The
        same effect can be produced if the code is
        compiled with the -Os option to the compiler."
}

cdl_component CYGPKG_LIBC_STRING_STRTOK {
    display       "strtok"
    flavor        none
    description   "
        These options control the behaviour of the
        strtok() and strtok_r() string tokenization
        functions."

    cdl_option CYGSEM_LIBC_PER_THREAD_STRTOK {
        display       "Per-thread strtok()"
        requires      CYGVAR_KERNEL_THREADS_DATA
        default_value 0
        description   "
            This option controls whether the string function
            strtok() has its state recorded on a per-thread
            basis rather than global. If this option is
            disabled, some per-thread space can be saved.
            Note there is also a POSIX-standard strtok_r()
            function to achieve a similar effect with user
            support. Enabling this option will use one slot
            of kernel per-thread data. You should ensure you
            have enough slots configured for all your
            per-thread data."
    }

    cdl_option CYGNUM_LIBC_STRTOK_TRACE_LEVEL {
        display       "Tracing level"
        flavor        data
        legal_values  0 to 1
        default_value 0
        description   "
            Trace verbosity level for debugging the <string.h>
            functions strtok() and strtok_r(). Increase this
            value to get additional trace output."
    }
}
