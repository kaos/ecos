# ====================================================================
#
#      hal_arm.cdl
#
#      ARM architectural HAL package configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      bartv
# Original data:  gthomas
# Contributors:
# Date:           1999-06-13
#
#####DESCRIPTIONEND####
#
# ====================================================================
cdl_package CYGPKG_HAL_ARM {
    display       "ARM architecture"
    parent        CYGPKG_HAL
    hardware
    include_dir   cyg/hal
    define_header hal_arm.h
    description   "
        The ARM architecture HAL package provides generic
        support for this processor architecture. It is also
        necessary to select a specific target platform HAL
        package."

    compile       hal_misc.c context.S arm_stub.c hal_syscall.c

    # The "-o file" is a workaround for CR100958 - without it the
    # output file would end up in the source directory under CygWin.
    # n.b. grep does not behave itself under win32
    make -priority 1 {
        arm.inc : <PACKAGE>/src/hal_mk_defs.c
        $(CC) $(CFLAGS) $(INCLUDE_PATH) -Wp,-MD,arm.tmp -o hal_mk_defs.tmp -S $<
        fgrep .equ hal_mk_defs.tmp | sed s/#// > $@
        @echo $@ ": \\" > $(notdir $@).deps
        @tail +2 arm.tmp >> $(notdir $@).deps
        @echo >> $(notdir $@).deps
        @rm arm.tmp hal_mk_defs.tmp
    }

    make {
        <PREFIX>/lib/vectors.o : <PACKAGE>/src/vectors.S
        $(CC) -Wp,-MD,vectors.tmp $(INCLUDE_PATH) $(CFLAGS) -c -o $@ $<
        @echo $@ ": \\" > $(notdir $@).deps
        @tail +2 vectors.tmp >> $(notdir $@).deps
        @echo >> $(notdir $@).deps
        @rm vectors.tmp
    }

    make {
        <PREFIX>/lib/target.ld: <PACKAGE>/src/arm.ld
        $(CC) -E -P -Wp,-MD,target.tmp -DEXTRAS=1 -xc $(INCLUDE_PATH) $(CFLAGS) -o $@ $<
        @echo $@ ": \\" > $(notdir $@).deps
        @tail +2 target.tmp >> $(notdir $@).deps
        @echo >> $(notdir $@).deps
        @rm target.tmp
    }

    cdl_interface CYGINT_HAL_ARM_THUMB_ARCH {
        display "The CPU architecture supports THUMB mode"
    }

    cdl_option CYGHWR_THUMB {
        display          "Enable Thumb instruction set"
        active_if        { CYGINT_HAL_ARM_THUMB_ARCH != 0 }
        default_value    0
        description      "
            Enable use of the Thumb instruction set."
    }

    # Note that when building a ROM monitor we include Thumb
    # interworking in order to support Thumb applications running
    # under a ARM ROM monitor.
    cdl_option CYGBLD_ARM_ENABLE_THUMB_INTERWORK {
        display       "Enable Thumb interworking compiler option"
        active_if        { CYGINT_HAL_ARM_THUMB_ARCH != 0 }
        default_value { (CYGHWR_THUMB || CYGSEM_HAL_ROM_MONITOR) }
        description "
            This option controls the use of -mthumb-interwork in the
            compiler flags. It defaults enabled in Thumb or ROM monitor
            configurations, but can be overridden for reduced memory
            footprint where interworking is not a requirement."
    }

    cdl_interface CYGINT_HAL_ARM_BIGENDIAN {
        display "The platform and architecture supports Big Endian operation"
    }

    cdl_option CYGHWR_HAL_ARM_BIGENDIAN {
        display          "Use big-endian mode"
        active_if        { CYGINT_HAL_ARM_BIGENDIAN != 0 }
        default_value    0
        description      "
            Use the CPU in big-endian mode."
    }

    cdl_interface CYGINT_HAL_ARM_ARCH_ARM7 {
        display "The platform uses a processor with an ARM7 core"
    }

    cdl_interface CYGINT_HAL_ARM_ARCH_ARM9 {
        display "The platform uses a processor with an ARM9 core"
    }

    cdl_interface CYGINT_HAL_ARM_ARCH_STRONGARM {
        display "The platform uses a processor with a StrongARM core"
    }

    cdl_interface CYGINT_HAL_ARM_ARCH_XSCALE {
        display "The platform uses a processor with a XScale core"
    }

    cdl_option CYGHWR_HAL_ARM_CPU_FAMILY {
        display       "ARM CPU family"
        flavor        data
        legal_values  { (CYGINT_HAL_ARM_ARCH_ARM7 != 0) ? "ARM7" : ""
                        (CYGINT_HAL_ARM_ARCH_ARM9 != 0) ? "ARM9" : ""
                        (CYGINT_HAL_ARM_ARCH_STRONGARM != 0) ? "StrongARM" : ""
                        (CYGINT_HAL_ARM_ARCH_XSCALE != 0) ? "XScale" : ""
                        "" }
        default_value  { (CYGINT_HAL_ARM_ARCH_ARM7 != 0) ? "ARM7" : 
                         (CYGINT_HAL_ARM_ARCH_ARM9 != 0) ? "ARM9" : 
                         (CYGINT_HAL_ARM_ARCH_STRONGARM != 0) ? "StrongARM" : 
                         (CYGINT_HAL_ARM_ARCH_XSCALE != 0) ? "XScale" :
                         "unknown" }
        no_define
        description   "
             It is possible to optimize code for different
             ARM CPU families. This option selects which CPU to
             optimize for on boards that support multiple CPU types."
    }

    cdl_option CYGHWR_HAL_ARM_DUMP_EXCEPTIONS {
        display          "Provide diagnostic dump for exceptions"
        requires         !CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
        default_value    0
        description      "
            Print messages about hardware exceptions, including
            raw exception frame dump and register contents."
    }

    cdl_option CYGIMP_HAL_PROCESS_ALL_EXCEPTIONS {
        display          "Process all exceptions with the eCos application"
        default_value    0
        description      "
           Normal RAM-based programs which do not include GDB stubs 
           defer processing of the illegal instruction exception to GDB.
           Setting this options allows the program to explicitly handle
           the illegal instruction exception itself.  Note: this will
           prevent the use of GDB to debug the application as breakpoints
           will no longer work."
    }

    cdl_option CYGBLD_LINKER_SCRIPT {
        display "Linker script"
        flavor data
	no_define
        calculated  { "src/arm.ld" }
    }

    cdl_interface CYGINT_HAL_ARM_MEM_REAL_REGION_TOP {
        display  "Implementations of hal_arm_mem_real_region_top()"
    }
}
