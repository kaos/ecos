# ====================================================================
#
#      wallclock_sh3.cdl
#
#      eCos wallclock SH3 RTC-module driver configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  nickg
# Contributors:
# Date:           2000-04-05
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVICES_WALLCLOCK_SH3 {
    parent        CYGPKG_IO_WALLCLOCK
    active_if     CYGPKG_IO_WALLCLOCK
    display       "SH3 RTC-module wallclock driver"
    requires      CYGPKG_HAL_SH
    hardware
    compile       wallclock_sh3.cxx
    define_proc {
        puts $::cdl_header "#undef CYGSEM_WALLCLOCK_SET_GET_MODE"
    }
    implements    CYGINT_WALLCLOCK_HW_IMPLEMENTATIONS
    active_if     CYGIMP_WALLCLOCK_HARDWARE

    cdl_option CYGIMP_WALLCLOCK_HARDWARE {
        parent    CYGPKG_IO_WALLCLOCK_IMPLEMENTATION
        display       "Hardware wallclock"
        default_value 1
        implements    CYGINT_WALLCLOCK_IMPLEMENTATIONS
    }

    cdl_component CYGPKG_DEVICES_WALLCLOCK_SH3_OPTIONS {
        display "SH3 RTC-module wallclock build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_DEVICES_WALLCLOCK_SH3_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the wallclock device. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_DEVICES_WALLCLOCK_SH3_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the wallclock device. These flags are removed from
                the set of global flags if present."
        }

    }
}
