# ====================================================================
#
#      ns_dp83902a_eth_drivers.cdl
#
#      Ethernet drivers - device support for NS DP83902A Ethernet
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000, 2001 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Contributors:   gthomas, jskov
# Date:           2001-06-13
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_NS_DP83902A {
    display       "NS DP83902A ethernet drivers"

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if     CYGPKG_IO_ETH_DRIVERS

    implements    CYGHWR_NET_DRIVERS

    active_if     CYGINT_DEVS_ETH_NS_DP83902A_REQUIRED

    include_dir   cyg/io
    description   "Ethernet driver for NS DP83902A (and DP8390) ethernet controller."
    compile       -library=libextras.a if_dp83902a.c

    define_proc {
        puts $::cdl_header "#include <pkgconf/system.h>";
        puts $::cdl_header "#include CYGDAT_DEVS_ETH_NS_DP83902A_CFG";
    }

    cdl_component CYGPKG_DEVS_ETH_DP83902A_OPTIONS {
        display "DP83902A ethernet driver build options"
        flavor  none
	no_define

        cdl_option CYGPKG_DEVS_ETH_DP83902A_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building the Cirrus Logic ethernet driver package.
                These flags are used in addition
                to the set of global flags."
        }
    }
}
