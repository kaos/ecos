# ====================================================================
#
#      time.cdl
#
#      C library time related configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  jlarmour
# Contributors:
# Date:           1999-07-06
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_option CYGSEM_LIBC_TIME_CLOCK_WORKING {
    display       "Working clock() function"
    requires      CYGFUN_KERNEL_THREADS_TIMER
    requires      CYGVAR_KERNEL_COUNTERS_CLOCK
    default_value 1
    description   "
        This option controls whether clock() will
        actually try and determine the process time
        usage. With this option disabled, clock() does
        not disappear, but will permanently return
        (clock_t)-1 as mandated by the ISO C standard."
}

cdl_option CYGSEM_LIBC_TIME_TIME_WORKING {
    display       "Working time() function"
    requires      CYGPKG_DEVICES_WALLCLOCK
    default_value 1
    description   "
        This option controls whether time() will
        actually try and determine the current calendar
        time. With this option disabled, time() does
        not disappear, but will permanently return
        (time_t)-1 as mandated by the ISO C standard."
}

cdl_option CYGSEM_LIBC_TIME_SETTIME_WORKING {
    display       "Working cyg_libc_time_settime() function"
    requires      CYGPKG_DEVICES_WALLCLOCK
    default_value 1
    description   "
        This option controls whether cyg_libc_time_settime()
        will actually try and set the current calendar
        time. With this option disabled,
        cyg_libc_time_settime() does not disappear, but
        will permanently return an error."
}

cdl_option CYGFUN_LIBC_TIME_POSIX {
    display       "POSIX time functions"
    default_value 1
    description   "
        Enabling this option allows the use of the
        following functions defined in POSIX 1003.1:
        asctime_r(), ctime_r(), gmtime_r(), and
        localtime_r()."
}

cdl_component CYGPKG_LIBC_TIME_ZONES {
    display       "Time zone offsets"
    flavor        none
    description   "
        These options control the default STandarD (STD)
        and Daylight Savings Time (DST)
        time offsets so that dates can be set correctly
        for the local environment."
    
    cdl_option CYGNUM_LIBC_TIME_DST_DEFAULT_STATE {
        display       "Default Daylight Savings Time state"
        flavor        data
        legal_values  -- -1 to 1
        default_value -- -1
        description   "
            This option controls whether the initial
            time environment is set up as STD, DST or
            unknown. Use the value 1 for DST, 0 for STD, 
            and (-1) for unknown. This can also be set at
            runtime using the cyg_libc_time_setdst()
            function."
    }

    cdl_option CYGNUM_LIBC_TIME_STD_DEFAULT_OFFSET {
        display       "Default Standard Time offset"
        flavor        data
        legal_values  -- -90000 to 90000
        default_value -- 0
        description   "
            This option controls the offset from UTC in
            seconds when in local Standard Time. This
            value can be positive or negative. It
            can also be set at run time using the
            cyg_libc_time_setzoneoffsets() function."
    }

    cdl_option CYGNUM_LIBC_TIME_DST_DEFAULT_OFFSET {
        display       "Default Daylight Savings Time offset"
        flavor        data
        legal_values  -- -90000 to 90000
        default_value -- 3600
        description   "
            This option controls the offset from UTC in
            seconds when in local Daylight Savings Time. This
            value can be positive or negative. It
            can also be set at run time using the
            cyg_libc_time_setzoneoffsets() function."
    }
}        

cdl_component CYGPKG_LIBC_TIME_INLINES {
    display       "Inline functions"
    flavor        none
    description   "
        These options control whether certain functions
        are available in inline form. This may lead to
        faster code at the expense of code space. But for
        some functions, or some functions with constant
        arguments, it may in fact lead to smaller code."

    cdl_option CYGIMP_LIBC_TIME_ASCTIME_INLINE {
        display       "asctime()"
        default_value 1
        description   "
            Allow the asctime() function to be inlined"
    }

    cdl_option CYGIMP_LIBC_TIME_CTIME_INLINE {
        display       "ctime()"
        default_value 1
        description   "
            Allow the ctime() function to be inlined"
    }

    cdl_option CYGIMP_LIBC_TIME_DIFFTIME_INLINE {
        display       "difftime()"
        default_value 1
        description   "
            Allow the difftime() function to be inlined"
    }

    cdl_option CYGIMP_LIBC_TIME_GMTIME_INLINE {
        display       "gmtime()"
        default_value 1
        description   "
            Allow the gmtime() function to be inlined"
    }

    cdl_option CYGIMP_LIBC_TIME_LOCALTIME_INLINE {
        display       "localtime()"
        default_value 1
        description   "
            Allow the localtime() function to be inlined"
    }

    cdl_option CYGIMP_LIBC_TIME_MKTIME_INLINE {
        display       "mktime()"
        default_value 1
        description   "
            Allow the mktime() function to be inlined"
    }

    cdl_option CYGIMP_LIBC_TIME_ASCTIME_R_INLINE {
        display       "asctime_r()"
        requires      CYGFUN_LIBC_TIME_POSIX
        default_value 1
        description   "
            Allow the asctime_r() function to be inlined"
    }

    cdl_option CYGIMP_LIBC_TIME_CTIME_R_INLINE {
        display       "ctime_r()"
        requires      CYGFUN_LIBC_TIME_POSIX
        default_value 1
        description   "
            Allow the ctime_r() function to be inlined"
    }

    cdl_option CYGIMP_LIBC_TIME_GMTIME_R_INLINE {
        display       "gmtime_r()"
        requires      CYGFUN_LIBC_TIME_POSIX
        default_value 1
        description   "
            Allow the gmtime_r() function to be inlined"
    }

    cdl_option CYGIMP_LIBC_TIME_LOCALTIME_R_INLINE {
        display       "localtime_r()"
        requires      CYGFUN_LIBC_TIME_POSIX
        default_value 1
        description   "
            Allow the localtime_r() function to be inlined"
    }
}
# FIXME: Also want "inline all" and "don't inline any" options which requires
# (or not) all the above, but
# if we do that then we will require the ones that also depend on
# CYGFUN_LIBC_TIME_POSIX :-( Wait for full CDL to fix this

cdl_option CYGNUM_LIBC_TIME_CLOCK_TRACE_LEVEL {
    display       "clock() tracing level"
    flavor        data
    legal_values  0 to 1
    default_value 0
    description   "
        Trace verbosity level for debugging the clock()
        function. Increase this value to get
        additional trace output when tracing is enabled."
}
