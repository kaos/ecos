# ====================================================================
#
#      usbs_serial.cdl
#
#      USB slave-side serial package.
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2008 Free Software Foundation, Inc.                        
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Frank M. Pagliughi (fmp), SoRo Systems, Inc.
# Contributors:
# Date:           2008-06-04
#
#####DESCRIPTIONEND####
# ====================================================================

cdl_package CYGPKG_IO_USB_SLAVE_SERIAL {
    display     "USB slave serial support"
    include_dir "cyg/io/usb"
    parent      CYGPKG_IO_USB_SLAVE
    requires    { CYGHWR_IO_USB_SLAVE_OUT_ENDPOINTS >= 1 }
    requires    { CYGHWR_IO_USB_SLAVE_IN_ENDPOINTS >= 1 }
    compile     usbs_serial.c
    implements  CYGINT_IO_USB_SLAVE_CLIENTS
#    doc         ref/io-usb-slave-eth.html
    
    description "
        The USB slave serial package supports the development of USB
        peripherals which mimic a serial connection to the host
        machine. Such a device creates a relatively simple upgrade to
        USB from a legacy serial connection, especially from the
        perspective of the host software and device drivers."

    cdl_option CYGDAT_IO_USB_SLAVE_CLASS_TYPE {
        display         "Serial USB Class"
        flavor          data
        default_value   { "ACM" }
        legal_values    { "ACM" "generic" }
        description     "
            The USB serial module can enumerate as either a generic
            (vendor-specific) usb device or a communications class ACM
            device. The generic device requires a pair of Bulk
            endpoints, while the ACM device also requires an Interrupt
            IN endpoint.  For a Windows host, the ACM configuration is
            required to use the standard 'usbser.sys' device driver,
            but for a Linux host, the generic configuration works, and
            saves the additional endpoint."
    }
    cdl_option CYGDAT_IO_USB_SLAVE_SERIAL_EP0 {
        display       "Name of EP0 structure"
        flavor        data               
        default_value { "usbs_at91_ep0" }
        description   "
            The name of the variable that contains the endpoint 0
            structure.  This should be set to the EP0 structure for
            the desired USB device driver such as usbs_at91_ep0,
            usbs_sa11x0_ep0, etc"
    }
    cdl_option CYGNUM_IO_USB_SLAVE_SERIAL_EP0_MAX_PACKET_SIZE {
        display       "The size of EP0"
        flavor        data
        default_value 8
        legal_values  { 8 16 64 } 
        description   "
            The size of the EP0 hardware buffer on the specific USB
            chip used."
    } 
    cdl_option CYGNUM_IO_USB_SLAVE_SERIAL_TX_EP_NUM {
        display       "Tx (USB IN) endpoint number"
        flavor        data
        default_value 1
        description   "
            The endpoint that should be used for the device-side
            transmitter, which is the USB IN direction."
    }
    cdl_option CYGDAT_IO_USB_SLAVE_SERIAL_TX_EP {
        display         "The Tx (USB IN) endpoint structure"
         flavor         data               
         default_value  { "usbs_at91_ep1" }
         description    "
             The endpoint structure that corresponds to the selected
             Tx endpoint number. This is dependent on the USBS device
             driver selected, and could be usbs_at91_ep1,
             usbs_sa11x0_ep1, etc"

    }
    cdl_option CYGNUM_IO_USB_SLAVE_SERIAL_RX_EP_NUM {
        display         "Rx (USB OUT) endpoint number"
        flavor          data
        default_value   2
        description     "
            The endpoint that should be used for the device-side
            receiver, which is the USB OUT direction."
    } 
    cdl_option CYGDAT_IO_USB_SLAVE_SERIAL_RX_EP {
        display         "The Rx (USB OUT) endpoint structure"
         flavor         data               
         default_value  { "usbs_at91_ep2" }
         description    "
             The endpoint structure that corresponds to the selected
             Rx endpoint number. This is dependent on the USBS device
             driver selected, and could be usbs_at91_ep2,
             usbs_sa11x0_ep2, etc"
    }
    cdl_option CYGNUM_IO_USB_SLAVE_SERIAL_INTR_EP_NUM {
        display         "Interrupt IN endpoint number"
        flavor          data
        default_value   3
        active_if       { CYGDAT_IO_USB_SLAVE_CLASS_TYPE == "ACM" }
        description     "
            The endpoint that should be used for the ACM Interrupt IN"
    }
    cdl_option CYGDAT_IO_USB_SLAVE_SERIAL_INTR_EP {
        display         "Interrupt IN endpoint structure"
         flavor         data               
         default_value  { "usbs_at91_ep3" }
         active_if      { CYGDAT_IO_USB_SLAVE_CLASS_TYPE == "ACM" }
         description    "
             The endpoint structure that corresponds to the selected ACM
             Interrupt IN endpoint."
    }
    cdl_option CYGNUM_IO_USB_SLAVE_SERIAL_VENDOR_ID {
        display       "USB Forum Vendor ID"
        flavor        data
        default_value 0xFFFF
        legal_values  1 to 0xFFFF
        description   "
            Each USB vendor has an Vendor ID allocated to it by the
            USB-IF organization.  Any arbitrary value can be selected
            for testing provided that it doesn't conflict with devices
            on the development host, but a device should NEVER be
            released publicly without a valid Vendor ID"

    }
    cdl_option CYGNUM_IO_USB_SLAVE_SERIAL_PRODUCT_ID {
        display       "USB product ID"
        flavor        data
        default_value 1
        legal_values  1 to 0xFFFF
        description   "
            You are free to select an arbitrary 16-bit Product ID for
            a device. The combination of Vendor ID and Product ID
            uniquely identified a USB device."
    }
    cdl_option CYGDAT_IO_USB_SLAVE_SERIAL_MFG_STR {
        display       "The Device Vendor's Name (Manufacturer String)"
        flavor        data
        default_value { "\"eCos\"" }
        description "
                The standard USB enumeration allows for a
                manufacturer's name which is normally reported to the
                user when the device is first plugged into the host."
    }
    cdl_option CYGDAT_IO_USB_SLAVE_SERIAL_PRODUCT_STR {
        display       "The Device Product Name"
        flavor        data
        default_value { "\"eCos USB Serial Device\"" }
        description "
                The standard USB enumeration allows for a product name
                which is normally reported to the user when the device
                is first plugged into the host."
    }

    cdl_option CYGOPT_IO_USB_SLAVE_SERIAL_BUSPOWERED {
        display       "The Device is bus powered"
        default_value 0
        flavor        bool
        description   "
            Tells the host whether the Device is a bus powered
            device or a self powered device."
    }
    cdl_option CYGNUM_IO_USB_SLAVE_SERIAL_CURRENTDRAW {
        display       "Maximum current (in mA) drawn from USB bus"
        flavor        data
        default_value 100
        legal_values  1 to 500
        requires      { (CYGNUM_IO_USB_SLAVE_SERIAL_CURRENTDRAW > 100) 
                         implies CYGOPT_IO_USB_SLAVE_SERIAL_BUSPOWERED }
        description   "
            The maximum current drawn by the Device from the USB bus.
            It should report the peak value. A self powered device
            can draw up to 100mA, a bus powered device can draw up to
            500mA. (If it is sometimes below 100mA and sometimes over,
            then a tranition could be done at runtime between self and
            bus powered modes, but that would be complicated and the
            device would have to return from configured to addressed
            state. For details, see the USB specification.)"
    }

    cdl_option  CYGBLD_IO_USB_SLAVE_SERIAL_DEBUG {
        display       "Enable debug output from the driver"
        default_value 0
        flavor        bool
        description   "
            The driver may produce debug output which can be
            useful to work out why it is not working as expected."
    }

    cdl_component CYGPKG_IO_USB_SLAVE_SERIAL_OPTIONS {
    display     "Build options"
    flavor      none

    description "
        Package-specific build options including control over compiler
        flags used only in building this package."

        cdl_option CYGPKG_IO_USB_SLAVE_SERIAL_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building this package. These flags are used in addition
                to the set of global flags."
        }
 
        cdl_option CYGPKG_IO_USB_SLAVE_SERIAL_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building this package. These flags are removed from
                the set of global flags if present."
        }
    

        cdl_component CYGBLD_IO_USB_SLAVE_SERIAL_EXAMPLES {
            display "Build example programs"
            no_define
            requires    { CYGPKG_IO_FILEIO }         
            requires    { CYGPKG_IO_SERIAL_DEVICES }         
            description "
                Enabling this option will cause the example programs
                to be built using the normal test case infrastructure.
                They are however not test cases and should not be used
                with any automatic test farm running all the
                tests. Hence this option is disabled by default."
            
             cdl_option CYGPKG_IO_USB_SLAVE_SERIAL_TESTS {
                 display "USBS serial example/test programs"
                 no_define
                 flavor data
                 calculated { "tests/usbserial_echo.c tests/usb2serial.c" }
                 description "
                     usbserial_echo will echo charactors received
                     over the usb serial port back to the sender.
                     usb2serial acts as a bridge between a USB serial
                     slave and a real serial port. It is hard coded to use
                     /dev/ser0."
             }
        }
    }
}
