# ====================================================================
#
#      flash_amd_am29f040b.cdl
#
#      FLASH memory - Hardware support for AMD AM29F040B
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Contributors:   gthomas, jskov
# Date:           2000-12-05
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_FLASH_AMD_AM29F040B {
    display       "AMD AM29F040B FLASH memory support"
    description   "FLASH memory device support for AMD AM29F040B"
    parent        CYGPKG_IO_FLASH
    active_if	  CYGPKG_IO_FLASH

    active_if     CYGINT_DEVS_FLASH_AMD_AM29F040B_REQUIRED

    implements    CYGHWR_IO_FLASH_DEVICE

    include_dir   .
    include_files ; # none _exported_ whatsoever

    compile       am29f040b_flash.c

    define_proc {
        puts $::cdl_header "#include <pkgconf/system.h>";
        puts $::cdl_header "#include CYGDAT_DEVS_FLASH_AMD_AM29F040B_CFG";
    }

    make -priority 1 {
        flash_query.o: $(REPOSITORY)/$(PACKAGE)/src/flash_query.c
        $(CC) -S $(INCLUDE_PATH) -mips2 -EB -fno-function-sections $(REPOSITORY)/$(PACKAGE)/src/flash_query.c
        echo "#include <cyg/io/plf_flash.inc>" > flash_query2.S
        cat  flash_query.s >> flash_query2.S
        echo "FUNC_END(flash_query_end)" >>flash_query2.S
        $(CC) -c $(INCLUDE_PATH) -mips2 -EB -G0 -o flash_query.o flash_query2.S
        $(AR) rcs $(PREFIX)/lib/libtarget.a flash_query.o
    }

    make -priority 1 {
        flash_erase_block.o: $(REPOSITORY)/$(PACKAGE)/src/flash_erase_block.c
        $(CC) -S $(INCLUDE_PATH) -mips2 -EB -fno-function-sections $(REPOSITORY)/$(PACKAGE)/src/flash_erase_block.c
        echo "#include <cyg/io/plf_flash.inc>" > flash_erase_block2.S
        cat  flash_erase_block.s >> flash_erase_block2.S
        echo "FUNC_END(flash_erase_block_end)" >>flash_erase_block2.S
        $(CC) -c $(INCLUDE_PATH) -mips2 -EB -G0 -o flash_erase_block.o flash_erase_block2.S
        $(AR) rcs $(PREFIX)/lib/libtarget.a flash_erase_block.o
    }

    make -priority 1 {
        flash_program_buf.o: $(REPOSITORY)/$(PACKAGE)/src/flash_program_buf.c
        $(CC) -S $(INCLUDE_PATH) -mips2 -EB -fno-function-sections $(REPOSITORY)/$(PACKAGE)/src/flash_program_buf.c
        echo "#include <cyg/io/plf_flash.inc>" > flash_program_buf2.S
        cat  flash_program_buf.s >> flash_program_buf2.S
        echo "FUNC_END(flash_program_buf_end)" >>flash_program_buf2.S
        $(CC) -c $(INCLUDE_PATH) -mips2 -EB -G0 -o flash_program_buf.o flash_program_buf2.S
        $(AR) rcs $(PREFIX)/lib/libtarget.a flash_program_buf.o
    }
}

