# ====================================================================
#
#      hal_powerpc_moab.cdl
#
#      PowerPC/MOAB board HAL package configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
## Copyright (C) 2002, 2003 Gary Thomas
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  hmt
# Contributors:   gthomas
# Date:           1999-11-02
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_POWERPC_MOAB {
    display       "TAMS MOAB (PowerPC 405GPr) board"
    parent        CYGPKG_HAL_POWERPC
    requires      CYGPKG_HAL_POWERPC_PPC40x
    define_header hal_powerpc_moab.h
    include_dir   cyg/hal
    description   "
        The MOAB HAL package provides the support needed to run
        eCos on a TAMS PowerPC 405GP board."

    compile       hal_aux.c moab.S

    implements    CYGINT_HAL_DEBUG_GDB_STUBS
    implements    CYGINT_HAL_DEBUG_GDB_STUBS_BREAK
    implements    CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT

    requires      CYGSEM_HAL_POWERPC_RESET_USES_JUMP        
    requires      { CYGHWR_HAL_POWERPC_PPC4XX == "405GP" }
# work around DCACHE problems - see errata for details, but
# basically, writethru mode is the only safe way to run this
    requires      { CYGSEM_HAL_DCACHE_STARTUP_MODE == "WRITETHRU" }
# having the MMU enabled just seems to cause no end of problems
    requires      { !CYGHWR_HAL_POWERPC_ENABLE_MMU }
#
    requires      { !CYGSEM_REDBOOT_FLASH_CONFIG || 
                    ((CYGHWR_REDBOOT_FLASH_CONFIG_MEDIA == "EEPROM") &&
                     (CYGNUM_REDBOOT_FLASH_CONFIG_SIZE == CYGNUM_HAL_EEPROM_SIZE) &&
                     (CYGNUM_REDBOOT_FLASH_STRING_SIZE == 64) &&
                     (CYGNUM_REDBOOT_FLASH_SCRIPT_SIZE == 256)) }
    requires      { !CYGPKG_REDBOOT || CYGBLD_REDBOOT_MAX_MEM_SEGMENTS == 2 }

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H   <pkgconf/hal_powerpc_ppc40x.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_powerpc_moab.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLF_IO_H   <cyg/hal/plf_io.h>"

	puts $::cdl_header "#define HAL_PLATFORM_CPU    \"PowerPC 405GPr\""
        puts $::cdl_header "#define HAL_PLATFORM_BOARD  \"TAMS MOAB\""
        puts $::cdl_header "#define HAL_PLATFORM_EXTRA  \"\""
    }

    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        legal_values  {"RAM" "ROM" "ROMRAM"}
        default_value {"RAM"}
	no_define
	define -file system.h CYG_HAL_STARTUP
        description   "
           This option is used to control where the application program will
           run, either from RAM or ROM (flash) memory.  ROM based applications
           must be self contained, while RAM applications will typically assume
           the existence of a debug environment, such as GDB stubs."
    }

    cdl_option CYGHWR_HAL_POWERPC_CPU_SPEED {
        display          "Development board clock speed (MHz)"
        flavor           data
        legal_values     250 333
        default_value    250
        description      "
           MOAB Development Boards have various system clock speeds
           depending on the processor and oscillator fitted.  Select 
           the clock speed appropriate for your board so that the system 
           can set the serial baud rate correctly, amongst other things."
   }

   cdl_option CYGHWR_HAL_POWERPC_MEM_SPEED {
        display          "Development board memory bus speed (MHz)"
        flavor           data
        legal_values     66
        default_value    66
        description      "
           MOAB Development Boards have various system clock speeds
           depending on the processor and oscillator fitted."
   }

    cdl_component CYGNUM_HAL_EEPROM_SIZE {
        display       "Size of EEPROM device"
        flavor        data
        legal_values  { 1024 2048 4096 }
        default_value { 2048 }
        description   "
           This option indicates the size (and type) of EEPROM fitted on the board"
    }

    cdl_component CYGSEM_HAL_IDE_SUPPORT {
        display       "HAL support for IDE disks"
        flavor        bool
        active_if     CYGPKG_IO_PCI
        default_value 1
        implements    CYGINT_HAL_PLF_IF_IDE
        compile       moab_ide.c
        description   "
           Enable this option to get support for IDE devices.  This is useful
           to allow RedBoot to boot directly from disk."
    }
    
    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        description   "
	    Global build options including control over
	    compiler flags, linker flags and choice of toolchain."


        parent  CYGPKG_NONE

        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "powerpc-eabi" }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { "-msoft-float -mcpu=405 -Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority" }
            description   "
                This option controls the global compiler flags which
                are used to compile all packages by
                default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { "-msoft-float -mcpu=405 -g -nostdlib -Wl,--gc-sections -Wl,-static" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }

        cdl_option CYGBLD_BUILD_GDB_STUBS {
            display "Build GDB stub ROM image"
            default_value 0
            requires { CYG_HAL_STARTUP == "ROM" }
            requires CYGSEM_HAL_ROM_MONITOR
            requires CYGBLD_BUILD_COMMON_GDB_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT
            requires CYGDBG_HAL_DEBUG_GDB_THREAD_SUPPORT
            requires ! CYGDBG_HAL_COMMON_INTERRUPTS_SAVE_MINIMUM_CONTEXT
            requires ! CYGDBG_HAL_COMMON_CONTEXT_SAVE_MINIMUM
            no_define
            description "
                This option enables the building of the GDB stubs for the
                board. The common HAL controls takes care of most of the
                build process, but the platform CDL takes care of creating
                an S-Record data file suitable for programming using
                the board's EPPC-Bug firmware monitor."

            make -priority 320 {
                <PREFIX>/bin/gdb_module.bin : <PREFIX>/bin/gdb_module.img
                $(OBJCOPY) -O srec --change-address=0x02000000 $< $(@:.bin=.srec)
                $(OBJCOPY) -O binary $< $@
            }
        }
    }

    cdl_component CYGPKG_HAL_POWERPC_MOAB_OPTIONS {
        display "MOAB build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_HAL_POWERPC_MOAB_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the MOAB HAL. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_HAL_POWERPC_MOAB_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the MOAB HAL. These flags are removed from
                the set of global flags if present."
        }

        cdl_option CYGPKG_HAL_POWERPC_MOAB_TESTS {
            display "MOAB tests"
            flavor  data
            no_define
            calculated { "tests/moabtime" }
            description   "
                This option specifies the set of tests for the MOAB HAL."
        }
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { CYG_HAL_STARTUP == "RAM" ? "powerpc_moab_ram" : \
                     CYG_HAL_STARTUP == "ROMRAM" ? "powerpc_moab_romram" : \
                                                "powerpc_moab_rom" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_powerpc_moab_ram.ldi>" : \
                         CYG_HAL_STARTUP == "ROMRAM" ? "<pkgconf/mlt_powerpc_moab_romram.ldi>" : \
                                                    "<pkgconf/mlt_powerpc_moab_rom.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_powerpc_moab_ram.h>" : \
                         CYG_HAL_STARTUP == "ROMRAM" ? "<pkgconf/mlt_powerpc_moab_romram.h>" : \
                                                    "<pkgconf/mlt_powerpc_moab_rom.h>" }
        }
    }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "ROM" || CYG_HAL_STARTUP == "ROMRAM" }
        description   "
            Enable this option if this program is to be used as a ROM monitor,
            i.e. applications will be loaded into RAM on the board, and this
            ROM monitor may process exceptions or interrupts generated from the
            application. This enables features such as utilizing a separate
            interrupt stack when exceptions are generated."
    }

    cdl_component CYGPKG_REDBOOT_HAL_OPTIONS {
        display       "Redboot HAL options"
        flavor        none
        no_define
        parent        CYGPKG_REDBOOT
        active_if     CYGPKG_REDBOOT
        description   "
            This option lists the target's requirements for a valid Redboot
            configuration."

        cdl_option CYGSEM_REDBOOT_PLF_LINUX_BOOT {
            active_if      CYGBLD_BUILD_REDBOOT_WITH_EXEC
            display        "Support booting Linux via RedBoot"
            flavor         bool
            default_value  1
            description    "
               This option enables RedBoot to support booting of a Linux kernel."

            compile plf_redboot_linux_exec.c
        }

        cdl_component CYGBLD_BUILD_REDBOOT_OBJS {
            display       "Build Redboot image(s)"
            active_if     CYGBLD_BUILD_REDBOOT
            default_value 1
            no_define
            description "This option enables the conversion of the Redboot ELF
                         image various formats which simplify further manipulatations.
                         The most basic of these forms is Motorola S-records, which
                         are simpler and more reliable than binary formats when used
                         for serial download."

            make -priority 325 {
                <PREFIX>/bin/redboot.srec : <PREFIX>/bin/redboot.elf
                $(OBJCOPY) -O srec $< $(@:.bin=.srec)
            }

            cdl_option CYGBLD_BUILD_REDBOOT_BIN {
                display       "Build RedBoot ROM/FLASH binary image"
                default_value { CYG_HAL_STARTUP != "RAM" }
                description "This option enables the conversion of the Redboot ELF
                             image to a binary image suitable for ROM/FLASH programming."
                make -priority 324 {
                    <PREFIX>/bin/redboot.bin : <PREFIX>/bin/redboot.elf
                    $(OBJCOPY) -O binary $< /tmp/__redboot.bin
                    make_MOAB_flash /tmp/__redboot.bin $@
                    rm -f /tmp/__redboot.bin
                }
            }
        }
    }
}
