# ====================================================================
#
#      flags.cdl
#
#      uITRON flags related configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  hmt
# Contributors:
# Date:           1999-07-07
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_option CYGNUM_UITRON_FLAGS {
    display       "Number of eventflags"
    flavor        data
    legal_values  1 to 65535
    default_value 5
    description   "
        The number of uITRON eventflag objects present in the system.
        Valid eventflag object IDs will range from 1 to this value."
}
cdl_component CYGPKG_UITRON_FLAGS_CREATE_DELETE {
    display       "Support create and delete"
    flavor        bool
    default_value 1
    description   "
        Support eventflag create and delete operations (cre_flg, del_flg).
        Otherwise all eventflags are created, up to the number specified above."

    cdl_option CYGNUM_UITRON_FLAGS_INITIALLY {
        display       "Number of eventflags created initially"
        flavor        data
        legal_values  0 to 65535
        default_value 5
        description   "
            The number of uITRON eventflags initially created.
            This number should not be more than the number
            of eventflags in the system, though setting it to a large
            value to mean 'all' is acceptable.
            Initially, only eventflags numbered 1 to this number exist;
            higher numbered ones must be created before use."
    }
}
